/***
* This code is a part of EvoApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under The MIT License.
* When used, please cite the following article(s): PRABAKARAN B. S., MRAZEK V., VASICEK Z., SEKANINA L., SHAFIQUE M. ApproxFPGAs: Embracing ASIC-based Approximate Arithmetic Components for FPGA-Based Systems. DAC 2020. 
***/
// MAE% = 0.036 %
// MAE = 24 
// WCE% = 0.13 %
// WCE = 83 
// WCRE% = 300.00 %
// EP% = 94.20 %
// MRE% = 1.19 %
// MSE = 885 
// FPGA_POWER = 1.1
// FPGA_DELAY = 9.7
// FPGA_LUT = 74

module mul8u_7G9 (
    A,
    B,
    O
);

input [7:0] A;
input [7:0] B;
output [15:0] O;

wire sig_21,sig_22,sig_23,sig_28,sig_29,sig_30,sig_31,sig_32,sig_36,sig_37,sig_38,sig_41,sig_43,sig_44,sig_45,sig_46,sig_47,sig_49,sig_50,sig_51;
wire sig_52,sig_53,sig_54,sig_55,sig_57,sig_58,sig_59,sig_60,sig_61,sig_62,sig_63,sig_64,sig_65,sig_66,sig_67,sig_68,sig_69,sig_70,sig_71,sig_72;
wire sig_73,sig_74,sig_75,sig_76,sig_77,sig_78,sig_79,sig_97,sig_98,sig_99,sig_100,sig_101,sig_102,sig_103,sig_104,sig_105,sig_106,sig_107,sig_108,sig_109;
wire sig_110,sig_111,sig_112,sig_113,sig_116,sig_117,sig_118,sig_121,sig_122,sig_123,sig_124,sig_125,sig_126,sig_127,sig_128,sig_129,sig_130,sig_131,sig_132,sig_133;
wire sig_134,sig_135,sig_136,sig_137,sig_138,sig_139,sig_140,sig_141,sig_142,sig_143,sig_144,sig_145,sig_146,sig_147,sig_150,sig_151,sig_162,sig_164,sig_165,sig_166;
wire sig_167,sig_168,sig_169,sig_170,sig_171,sig_172,sig_173,sig_174,sig_175,sig_176,sig_177,sig_178,sig_179,sig_180,sig_182,sig_183,sig_184,sig_185,sig_186,sig_187;
wire sig_188,sig_189,sig_190,sig_191,sig_192,sig_193,sig_194,sig_195,sig_196,sig_197,sig_198,sig_199,sig_200,sig_201,sig_202,sig_203,sig_204,sig_205,sig_206,sig_207;
wire sig_208,sig_209,sig_210,sig_211,sig_212,sig_213,sig_214,sig_215,sig_216,sig_217,sig_218,sig_228,sig_229,sig_230,sig_231,sig_232,sig_233,sig_234,sig_235,sig_236;
wire sig_237,sig_238,sig_239,sig_240,sig_241,sig_242,sig_243,sig_244,sig_245,sig_246,sig_247,sig_248,sig_249,sig_250,sig_251,sig_252,sig_253,sig_254,sig_255,sig_256;
wire sig_263,sig_264,sig_265,sig_266,sig_267,sig_268,sig_269,sig_270,sig_271,sig_272,sig_273,sig_274,sig_275,sig_276,sig_277,sig_278,sig_279,sig_280,sig_281,sig_282;
wire sig_283,sig_284,sig_285,sig_286,sig_287,sig_288,sig_289,sig_290,sig_291,sig_292,sig_293,sig_294,sig_295,sig_296,sig_297,sig_298,sig_299,sig_328,sig_329,sig_330;
wire sig_331,sig_332,sig_333,sig_334,sig_335,sig_336,sig_337,sig_338,sig_339,sig_340,sig_341,sig_342,sig_343,sig_344,sig_384,sig_385,sig_386,sig_387,sig_388,sig_389;
wire sig_390,sig_391,sig_392,sig_393,sig_394,sig_395,sig_397,sig_398,sig_400,sig_401,sig_404,sig_405,sig_406,sig_407,sig_409,sig_410,sig_415,sig_416,sig_417,sig_418;
wire sig_419,sig_420,sig_421,sig_423,sig_424,sig_425,sig_428,sig_429;

assign sig_21 = B[5] & A[0];
assign sig_22 = B[6] & A[0];
assign sig_23 = B[7] & A[0];
assign sig_28 = B[4] & A[1];
assign sig_29 = B[5] & A[1];
assign sig_30 = B[6] & A[1];
assign sig_31 = B[7] & A[1];
assign sig_32 = B[2] & A[3];
assign sig_36 = B[4] & A[2];
assign sig_37 = B[5] & A[2];
assign sig_38 = B[6] & A[2];
assign sig_41 = B[3] & A[2];
assign sig_43 = B[3] & A[3];
assign sig_44 = B[4] & A[3];
assign sig_45 = B[5] & A[3];
assign sig_46 = B[6] & A[3];
assign sig_47 = B[7] & A[3];
assign sig_49 = B[1] & A[4];
assign sig_50 = B[2] & A[4];
assign sig_51 = B[3] & A[4];
assign sig_52 = B[4] & A[4];
assign sig_53 = B[5] & A[4];
assign sig_54 = B[6] & A[4];
assign sig_55 = B[7] & A[4];
assign sig_57 = B[1] & A[5];
assign sig_58 = B[2] & A[5];
assign sig_59 = B[3] & A[5];
assign sig_60 = B[4] & A[5];
assign sig_61 = B[5] & A[5];
assign sig_62 = B[6] & A[5];
assign sig_63 = B[7] & A[5];
assign sig_64 = B[0] & A[6];
assign sig_65 = B[1] & A[6];
assign sig_66 = B[2] & A[6];
assign sig_67 = B[3] & A[6];
assign sig_68 = B[4] & A[6];
assign sig_69 = B[5] & A[6];
assign sig_70 = B[6] & A[6];
assign sig_71 = B[7] & A[6];
assign sig_72 = B[0] & A[7];
assign sig_73 = B[1] & A[7];
assign sig_74 = B[2] & A[7];
assign sig_75 = B[3] & A[7];
assign sig_76 = B[4] & A[7];
assign sig_77 = B[5] & A[7];
assign sig_78 = B[6] & A[7];
assign sig_79 = B[7] & A[7];
assign sig_97 = sig_21 | sig_28;
assign sig_98 = sig_21 & sig_28;
assign sig_99 = sig_97 & sig_41;
assign sig_100 = sig_97 | sig_41;
assign sig_101 = sig_98 | sig_99;
assign sig_102 = sig_22 ^ sig_29;
assign sig_103 = sig_22 & sig_29;
assign sig_104 = sig_102 & sig_36;
assign sig_105 = sig_102 ^ sig_36;
assign sig_106 = sig_103 | sig_104;
assign sig_107 = sig_23 ^ sig_30;
assign sig_108 = sig_23 & sig_30;
assign sig_109 = sig_107 & sig_37;
assign sig_110 = sig_107 ^ sig_37;
assign sig_111 = sig_108 | sig_109;
assign sig_112 = sig_31 & sig_38;
assign sig_113 = sig_31 ^ sig_38;
assign sig_116 = sig_32 | sig_49;
assign sig_117 = sig_32 & sig_49;
assign sig_118 = sig_116 & B[0];
assign sig_121 = sig_43 ^ sig_50;
assign sig_122 = sig_43 & sig_50;
assign sig_123 = sig_121 & sig_57;
assign sig_124 = sig_121 ^ sig_57;
assign sig_125 = sig_122 | sig_123;
assign sig_126 = sig_44 ^ sig_51;
assign sig_127 = sig_44 & sig_51;
assign sig_128 = sig_126 & sig_58;
assign sig_129 = sig_126 ^ sig_58;
assign sig_130 = sig_127 | sig_128;
assign sig_131 = sig_45 ^ sig_52;
assign sig_132 = sig_45 & sig_52;
assign sig_133 = sig_131 & sig_59;
assign sig_134 = sig_131 ^ sig_59;
assign sig_135 = sig_132 | sig_133;
assign sig_136 = sig_46 ^ sig_53;
assign sig_137 = sig_46 & sig_53;
assign sig_138 = sig_136 & sig_60;
assign sig_139 = sig_136 ^ sig_60;
assign sig_140 = sig_137 | sig_138;
assign sig_141 = sig_47 ^ sig_54;
assign sig_142 = sig_47 & sig_54;
assign sig_143 = sig_141 & sig_61;
assign sig_144 = sig_141 ^ sig_61;
assign sig_145 = sig_142 | sig_143;
assign sig_146 = sig_55 & sig_62;
assign sig_147 = sig_55 ^ sig_62;
assign sig_150 = sig_105 | sig_101;
assign sig_151 = B[7] & A[2];
assign sig_162 = A[3] & B[1];
assign sig_164 = sig_100 | sig_162;
assign sig_165 = sig_105 ^ sig_101;
assign sig_166 = sig_105 & sig_101;
assign sig_167 = sig_150 & sig_124;
assign sig_168 = sig_165 ^ sig_124;
assign sig_169 = sig_166 | sig_167;
assign sig_170 = sig_110 ^ sig_106;
assign sig_171 = sig_110 & sig_106;
assign sig_172 = sig_170 & sig_129;
assign sig_173 = sig_170 ^ sig_129;
assign sig_174 = sig_171 | sig_172;
assign sig_175 = sig_113 ^ sig_111;
assign sig_176 = sig_113 & sig_111;
assign sig_177 = sig_175 & sig_134;
assign sig_178 = sig_175 ^ sig_134;
assign sig_179 = sig_176 | sig_177;
assign sig_180 = sig_151 ^ sig_112;
assign sig_182 = sig_151 & sig_139;
assign sig_183 = sig_180 ^ sig_139;
assign sig_184 = sig_112 | sig_182;
assign sig_185 = sig_118 ^ sig_64;
assign sig_186 = sig_118 & A[6];
assign sig_187 = sig_125 ^ sig_65;
assign sig_188 = sig_125 & sig_65;
assign sig_189 = sig_187 & sig_72;
assign sig_190 = sig_187 ^ sig_72;
assign sig_191 = sig_188 | sig_189;
assign sig_192 = sig_130 ^ sig_66;
assign sig_193 = sig_130 & sig_66;
assign sig_194 = sig_192 & sig_73;
assign sig_195 = sig_192 ^ sig_73;
assign sig_196 = sig_193 | sig_194;
assign sig_197 = sig_135 ^ sig_67;
assign sig_198 = sig_135 & sig_67;
assign sig_199 = sig_197 & sig_74;
assign sig_200 = sig_197 ^ sig_74;
assign sig_201 = sig_198 | sig_199;
assign sig_202 = sig_140 ^ sig_68;
assign sig_203 = sig_140 & sig_68;
assign sig_204 = sig_202 & sig_75;
assign sig_205 = sig_202 ^ sig_75;
assign sig_206 = sig_203 | sig_204;
assign sig_207 = sig_145 ^ sig_69;
assign sig_208 = sig_145 & sig_69;
assign sig_209 = sig_207 & sig_76;
assign sig_210 = sig_207 ^ sig_76;
assign sig_211 = sig_208 | sig_209;
assign sig_212 = sig_146 ^ sig_70;
assign sig_213 = sig_146 & A[6];
assign sig_214 = sig_212 & sig_77;
assign sig_215 = sig_212 ^ sig_77;
assign sig_216 = sig_213 | sig_214;
assign sig_217 = sig_71 & B[6];
assign sig_218 = sig_71 ^ sig_78;
assign sig_228 = sig_168 ^ sig_164;
assign sig_229 = sig_168 & sig_164;
assign sig_230 = sig_228 & sig_185;
assign sig_231 = sig_228 ^ sig_185;
assign sig_232 = sig_229 | sig_230;
assign sig_233 = sig_173 ^ sig_169;
assign sig_234 = sig_173 & sig_169;
assign sig_235 = sig_233 & sig_190;
assign sig_236 = sig_233 ^ sig_190;
assign sig_237 = sig_234 | sig_235;
assign sig_238 = sig_178 ^ sig_174;
assign sig_239 = sig_178 & sig_174;
assign sig_240 = sig_238 & sig_195;
assign sig_241 = sig_238 ^ sig_195;
assign sig_242 = sig_239 | sig_240;
assign sig_243 = sig_183 ^ sig_179;
assign sig_244 = sig_183 & sig_179;
assign sig_245 = sig_243 & sig_200;
assign sig_246 = sig_243 ^ sig_200;
assign sig_247 = sig_244 | sig_245;
assign sig_248 = sig_144 ^ sig_184;
assign sig_249 = sig_144 & sig_184;
assign sig_250 = sig_248 & sig_205;
assign sig_251 = sig_248 ^ sig_205;
assign sig_252 = sig_249 | sig_250;
assign sig_253 = sig_147 & sig_210;
assign sig_254 = sig_147 ^ sig_210;
assign sig_255 = sig_63 & sig_215;
assign sig_256 = sig_63 ^ sig_215;
assign sig_263 = sig_236 ^ sig_232;
assign sig_264 = sig_236 & sig_232;
assign sig_265 = sig_263 & sig_186;
assign sig_266 = sig_263 ^ sig_186;
assign sig_267 = sig_264 | sig_265;
assign sig_268 = sig_241 ^ sig_237;
assign sig_269 = sig_241 & sig_237;
assign sig_270 = sig_268 & sig_191;
assign sig_271 = sig_268 ^ sig_191;
assign sig_272 = sig_269 | sig_270;
assign sig_273 = sig_246 ^ sig_242;
assign sig_274 = sig_246 & sig_242;
assign sig_275 = sig_273 & sig_196;
assign sig_276 = sig_273 ^ sig_196;
assign sig_277 = sig_274 | sig_275;
assign sig_278 = sig_251 ^ sig_247;
assign sig_279 = sig_251 & sig_247;
assign sig_280 = sig_278 & sig_201;
assign sig_281 = sig_278 ^ sig_201;
assign sig_282 = sig_279 | sig_280;
assign sig_283 = sig_254 ^ sig_252;
assign sig_284 = sig_254 & sig_252;
assign sig_285 = sig_283 & sig_206;
assign sig_286 = sig_283 ^ sig_206;
assign sig_287 = sig_284 | sig_285;
assign sig_288 = sig_256 ^ sig_253;
assign sig_289 = sig_256 & sig_253;
assign sig_290 = sig_288 & sig_211;
assign sig_291 = sig_288 ^ sig_211;
assign sig_292 = sig_289 | sig_290;
assign sig_293 = sig_218 ^ sig_255;
assign sig_294 = sig_218 & sig_255;
assign sig_295 = sig_293 & sig_216;
assign sig_296 = sig_293 ^ sig_216;
assign sig_297 = sig_294 | sig_295;
assign sig_298 = A[7] & sig_217;
assign sig_299 = sig_79 ^ sig_298;
assign sig_328 = sig_271 ^ sig_267;
assign sig_329 = sig_271 & sig_267;
assign sig_330 = sig_276 ^ sig_272;
assign sig_331 = sig_276 & sig_272;
assign sig_332 = sig_330 & sig_329;
assign sig_333 = sig_330 ^ sig_329;
assign sig_334 = sig_331 | sig_332;
assign sig_335 = sig_281 ^ sig_277;
assign sig_336 = sig_281 & sig_277;
assign sig_337 = sig_335 & sig_334;
assign sig_338 = sig_335 ^ sig_334;
assign sig_339 = sig_336 | sig_337;
assign sig_340 = sig_286 ^ sig_282;
assign sig_341 = sig_286 & sig_282;
assign sig_342 = sig_340 & sig_339;
assign sig_343 = sig_340 ^ sig_339;
assign sig_344 = sig_341 | sig_342;
assign sig_384 = ~sig_344;
assign sig_385 = sig_291 & sig_287;
assign sig_386 = sig_296 ^ sig_292;
assign sig_387 = sig_296 & sig_292;
assign sig_388 = sig_386 & sig_385;
assign sig_389 = sig_386 ^ sig_385;
assign sig_390 = sig_387 | sig_388;
assign sig_391 = sig_299 ^ sig_297;
assign sig_392 = sig_299 & sig_297;
assign sig_393 = sig_391 & sig_390;
assign sig_394 = sig_391 ^ sig_390;
assign sig_395 = sig_392 | sig_393;
assign sig_397 = sig_298 | sig_395;
assign sig_398 = sig_291 ^ sig_287;
assign sig_400 = ~sig_398;
assign sig_401 = sig_385 | sig_398;
assign sig_404 = sig_386 & sig_401;
assign sig_405 = sig_386 ^ sig_401;
assign sig_406 = sig_390 | sig_404;
assign sig_407 = ~sig_344;
assign sig_409 = sig_391 & sig_406;
assign sig_410 = sig_391 ^ sig_406;
assign sig_415 = sig_398 & sig_407;
assign sig_416 = sig_400 & sig_344;
assign sig_417 = sig_415 | sig_416;
assign sig_418 = ~sig_344;
assign sig_419 = sig_389 & sig_418;
assign sig_420 = sig_405 & sig_344;
assign sig_421 = sig_419 | sig_420;
assign sig_423 = sig_394 & sig_384;
assign sig_424 = sig_410 & sig_344;
assign sig_425 = sig_423 | sig_424;
assign sig_428 = sig_409 & sig_344;
assign sig_429 = sig_397 | sig_428;

assign O[15] = sig_429;
assign O[14] = sig_425;
assign O[13] = sig_421;
assign O[12] = sig_417;
assign O[11] = sig_343;
assign O[10] = sig_338;
assign O[9] = sig_333;
assign O[8] = sig_328;
assign O[7] = sig_266;
assign O[6] = sig_231;
assign O[5] = sig_117;
assign O[4] = sig_29;
assign O[3] = sig_50;
assign O[2] = sig_106;
assign O[1] = sig_201;
assign O[0] = sig_395;

endmodule


