/***
* This code is a part of EvoApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under The MIT License.
* When used, please cite the following article(s): PRABAKARAN B. S., MRAZEK V., VASICEK Z., SEKANINA L., SHAFIQUE M. ApproxFPGAs: Embracing ASIC-based Approximate Arithmetic Components for FPGA-Based Systems. DAC 2020. 
***/
// MAE% = 1.95 %
// MAE = 83853312 
// WCE% = 7.81 %
// WCE = 335413249 
// WCRE% = 100.00 %
// EP% = 100.00 %
// MRE% = 19.30 %
// MSE = 10697.458e12 
// FPGA_POWER = 0.41
// FPGA_DELAY = 9.1
// FPGA_LUT = 17


module mul16u_GRC ( A, B, O );
  input [15:0] A;
  input [15:0] B;
  output [31:0] O;

  wire C_13_11,C_13_12,C_13_13,C_13_14,C_14_10,C_14_11,C_14_12,C_14_13,C_14_14,C_15_10,C_15_11,C_15_12,C_15_13,C_15_14,C_15_9,S_12_12,S_12_13,S_12_14,S_12_15,S_13_11,S_13_12,S_13_13,S_13_14,S_13_15,S_14_10,S_14_11,S_14_12,S_14_13,S_14_14,S_14_15,S_15_10,S_15_11,S_15_12,S_15_13,S_15_14,S_15_15,S_15_9,S_16_10,S_16_11,S_16_12,S_16_13,S_16_14,S_16_15,S_16_8,S_16_9;

  assign S_12_12 = (A[12] & B[12]);
  assign S_12_13 = (A[12] & B[13]);
  assign S_12_14 = (A[12] & B[14]);
  assign S_12_15 = (A[12] & B[15]);
  HAX1 U497940 (.A(S_12_12), .B((A[13] & B[11])), .YS(S_13_11), .YC(C_13_11));
  HAX1 U497941 (.A(S_12_13), .B((A[13] & B[12])), .YS(S_13_12), .YC(C_13_12));
  HAX1 U497942 (.A(S_12_14), .B((A[13] & B[13])), .YS(S_13_13), .YC(C_13_13));
  HAX1 U497943 (.A(S_12_15), .B((A[13] & B[14])), .YS(S_13_14), .YC(C_13_14));
  assign S_13_15 = (A[13] & B[15]);
  HAX1 U497955 (.A(S_13_11), .B((A[14] & B[10])), .YS(S_14_10), .YC(C_14_10));
  FAX1 U497956 (.A(S_13_12), .B(C_13_11), .C((A[14] & B[11])), .YS(S_14_11), .YC(C_14_11));
  FAX1 U497957 (.A(S_13_13), .B(C_13_12), .C((A[14] & B[12])), .YS(S_14_12), .YC(C_14_12));
  FAX1 U497958 (.A(S_13_14), .B(C_13_13), .C((A[14] & B[13])), .YS(S_14_13), .YC(C_14_13));
  FAX1 U497959 (.A(S_13_15), .B(C_13_14), .C((A[14] & B[14])), .YS(S_14_14), .YC(C_14_14));
  assign S_14_15 = (A[14] & B[15]);
  HAX1 U497970 (.A(S_14_10), .B((A[15] & B[9])), .YS(S_15_9), .YC(C_15_9));
  FAX1 U497971 (.A(S_14_11), .B(C_14_10), .C((A[15] & B[10])), .YS(S_15_10), .YC(C_15_10));
  FAX1 U497972 (.A(S_14_12), .B(C_14_11), .C((A[15] & B[11])), .YS(S_15_11), .YC(C_15_11));
  FAX1 U497973 (.A(S_14_13), .B(C_14_12), .C((A[15] & B[12])), .YS(S_15_12), .YC(C_15_12));
  FAX1 U497974 (.A(S_14_14), .B(C_14_13), .C((A[15] & B[13])), .YS(S_15_13), .YC(C_15_13));
  FAX1 U497975 (.A(S_14_15), .B(C_14_14), .C((A[15] & B[14])), .YS(S_15_14), .YC(C_15_14));
  assign S_15_15 = (A[15] & B[15]);
  assign {S_16_15, S_16_14, S_16_13, S_16_12, S_16_11, S_16_10, S_16_9, S_16_8} = {C_15_14, C_15_13, C_15_12, C_15_11, C_15_10, C_15_9, 1'b0} + {S_15_15, S_15_14, S_15_13, S_15_12, S_15_11, S_15_10, S_15_9};
  assign O = {S_16_15,S_16_14,S_16_13,S_16_12,S_16_11,S_16_10,S_16_9,S_16_8,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};

endmodule

