/***
* This code is a part of EvoApproxLib library (ehw.fit.vutbr.cz/approxlib) distributed under The MIT License.
* When used, please cite the following article(s): PRABAKARAN B. S., MRAZEK V., VASICEK Z., SEKANINA L., SHAFIQUE M. ApproxFPGAs: Embracing ASIC-based Approximate Arithmetic Components for FPGA-Based Systems. DAC 2020. 
***/
// MAE% = 0.000061 %
// MAE = 2606 
// WCE% = 0.00039 %
// WCE = 16653 
// WCRE% = 3100.00 %
// EP% = 99.93 %
// MRE% = 0.0044 %
// MSE = 11039.017e3 
// FPGA_POWER = 6.9
// FPGA_DELAY = 15
// FPGA_LUT = 349

module mul16u_01G (
	A,
	B,
	Z
);

input [15:0] A;
input [15:0] B;
output [31:0] Z;

wire sig_32;
wire sig_33;
wire sig_34;
wire sig_36;
wire sig_37;
wire sig_38;
wire sig_39;
wire sig_40;
wire sig_41;
wire sig_42;
wire sig_43;
wire sig_44;
wire sig_45;
wire sig_46;
wire sig_47;
wire sig_49;
wire sig_50;
wire sig_52;
wire sig_54;
wire sig_55;
wire sig_56;
wire sig_57;
wire sig_58;
wire sig_59;
wire sig_60;
wire sig_62;
wire sig_64;
wire sig_66;
wire sig_67;
wire sig_69;
wire sig_70;
wire sig_71;
wire sig_72;
wire sig_73;
wire sig_74;
wire sig_75;
wire sig_76;
wire sig_77;
wire sig_78;
wire sig_79;
wire sig_80;
wire sig_84;
wire sig_85;
wire sig_86;
wire sig_87;
wire sig_88;
wire sig_90;
wire sig_91;
wire sig_92;
wire sig_93;
wire sig_94;
wire sig_95;
wire sig_96;
wire sig_97;
wire sig_98;
wire sig_99;
wire sig_100;
wire sig_101;
wire sig_102;
wire sig_103;
wire sig_104;
wire sig_105;
wire sig_107;
wire sig_108;
wire sig_109;
wire sig_110;
wire sig_111;
wire sig_112;
wire sig_115;
wire sig_117;
wire sig_119;
wire sig_120;
wire sig_123;
wire sig_124;
wire sig_125;
wire sig_126;
wire sig_127;
wire sig_128;
wire sig_129;
wire sig_131;
wire sig_132;
wire sig_133;
wire sig_134;
wire sig_137;
wire sig_138;
wire sig_140;
wire sig_141;
wire sig_142;
wire sig_143;
wire sig_145;
wire sig_146;
wire sig_147;
wire sig_148;
wire sig_149;
wire sig_150;
wire sig_151;
wire sig_152;
wire sig_153;
wire sig_154;
wire sig_155;
wire sig_157;
wire sig_158;
wire sig_160;
wire sig_161;
wire sig_162;
wire sig_163;
wire sig_164;
wire sig_168;
wire sig_169;
wire sig_170;
wire sig_171;
wire sig_173;
wire sig_174;
wire sig_176;
wire sig_177;
wire sig_179;
wire sig_180;
wire sig_181;
wire sig_182;
wire sig_183;
wire sig_186;
wire sig_187;
wire sig_188;
wire sig_189;
wire sig_191;
wire sig_194;
wire sig_195;
wire sig_196;
wire sig_197;
wire sig_198;
wire sig_201;
wire sig_203;
wire sig_206;
wire sig_208;
wire sig_210;
wire sig_211;
wire sig_212;
wire sig_213;
wire sig_214;
wire sig_215;
wire sig_217;
wire sig_218;
wire sig_219;
wire sig_220;
wire sig_223;
wire sig_224;
wire sig_225;
wire sig_226;
wire sig_229;
wire sig_230;
wire sig_233;
wire sig_234;
wire sig_235;
wire sig_236;
wire sig_239;
wire sig_240;
wire sig_244;
wire sig_245;
wire sig_246;
wire sig_247;
wire sig_248;
wire sig_249;
wire sig_250;
wire sig_252;
wire sig_253;
wire sig_254;
wire sig_256;
wire sig_257;
wire sig_259;
wire sig_260;
wire sig_261;
wire sig_263;
wire sig_264;
wire sig_266;
wire sig_269;
wire sig_270;
wire sig_271;
wire sig_272;
wire sig_273;
wire sig_274;
wire sig_276;
wire sig_278;
wire sig_279;
wire sig_281;
wire sig_283;
wire sig_284;
wire sig_285;
wire sig_286;
wire sig_287;
wire sig_288;
wire sig_290;
wire sig_291;
wire sig_292;
wire sig_295;
wire sig_297;
wire sig_299;
wire sig_300;
wire sig_301;
wire sig_302;
wire sig_303;
wire sig_304;
wire sig_305;
wire sig_306;
wire sig_308;
wire sig_309;
wire sig_311;
wire sig_312;
wire sig_315;
wire sig_316;
wire sig_317;
wire sig_318;
wire sig_319;
wire sig_320;
wire sig_321;
wire sig_324;
wire sig_326;
wire sig_328;
wire sig_329;
wire sig_330;
wire sig_331;
wire sig_332;
wire sig_333;
wire sig_334;
wire sig_335;
wire sig_336;
wire sig_337;
wire sig_338;
wire sig_339;
wire sig_340;
wire sig_341;
wire sig_343;
wire sig_345;
wire sig_346;
wire sig_347;
wire sig_348;
wire sig_349;
wire sig_351;
wire sig_352;
wire sig_353;
wire sig_354;
wire sig_355;
wire sig_356;
wire sig_359;
wire sig_360;
wire sig_361;
wire sig_364;
wire sig_365;
wire sig_366;
wire sig_367;
wire sig_368;
wire sig_369;
wire sig_371;
wire sig_372;
wire sig_373;
wire sig_374;
wire sig_375;
wire sig_376;
wire sig_378;
wire sig_379;
wire sig_380;
wire sig_381;
wire sig_382;
wire sig_383;
wire sig_384;
wire sig_385;
wire sig_388;
wire sig_390;
wire sig_391;
wire sig_393;
wire sig_394;
wire sig_395;
wire sig_396;
wire sig_397;
wire sig_398;
wire sig_401;
wire sig_402;
wire sig_403;
wire sig_404;
wire sig_405;
wire sig_406;
wire sig_407;
wire sig_408;
wire sig_410;
wire sig_413;
wire sig_414;
wire sig_415;
wire sig_417;
wire sig_419;
wire sig_420;
wire sig_421;
wire sig_422;
wire sig_423;
wire sig_426;
wire sig_427;
wire sig_428;
wire sig_429;
wire sig_430;
wire sig_432;
wire sig_433;
wire sig_434;
wire sig_437;
wire sig_438;
wire sig_439;
wire sig_440;
wire sig_442;
wire sig_443;
wire sig_444;
wire sig_446;
wire sig_447;
wire sig_448;
wire sig_449;
wire sig_451;
wire sig_453;
wire sig_454;
wire sig_458;
wire sig_460;
wire sig_461;
wire sig_462;
wire sig_463;
wire sig_466;
wire sig_467;
wire sig_468;
wire sig_469;
wire sig_470;
wire sig_472;
wire sig_473;
wire sig_474;
wire sig_475;
wire sig_476;
wire sig_477;
wire sig_481;
wire sig_482;
wire sig_485;
wire sig_486;
wire sig_487;
wire sig_488;
wire sig_489;
wire sig_490;
wire sig_491;
wire sig_492;
wire sig_493;
wire sig_494;
wire sig_495;
wire sig_496;
wire sig_497;
wire sig_498;
wire sig_500;
wire sig_501;
wire sig_502;
wire sig_503;
wire sig_504;
wire sig_505;
wire sig_506;
wire sig_507;
wire sig_508;
wire sig_509;
wire sig_510;
wire sig_511;
wire sig_512;
wire sig_513;
wire sig_514;
wire sig_515;
wire sig_516;
wire sig_517;
wire sig_518;
wire sig_519;
wire sig_520;
wire sig_521;
wire sig_522;
wire sig_523;
wire sig_524;
wire sig_525;
wire sig_526;
wire sig_527;
wire sig_529;
wire sig_530;
wire sig_532;
wire sig_533;
wire sig_534;
wire sig_535;
wire sig_536;
wire sig_537;
wire sig_538;
wire sig_539;
wire sig_540;
wire sig_541;
wire sig_542;
wire sig_544;
wire sig_545;
wire sig_546;
wire sig_548;
wire sig_549;
wire sig_550;
wire sig_551;
wire sig_552;
wire sig_553;
wire sig_554;
wire sig_555;
wire sig_556;
wire sig_557;
wire sig_558;
wire sig_559;
wire sig_560;
wire sig_561;
wire sig_563;
wire sig_564;
wire sig_565;
wire sig_567;
wire sig_568;
wire sig_570;
wire sig_571;
wire sig_572;
wire sig_573;
wire sig_574;
wire sig_577;
wire sig_578;
wire sig_579;
wire sig_580;
wire sig_581;
wire sig_582;
wire sig_585;
wire sig_586;
wire sig_587;
wire sig_588;
wire sig_589;
wire sig_590;
wire sig_592;
wire sig_594;
wire sig_595;
wire sig_596;
wire sig_597;
wire sig_598;
wire sig_599;
wire sig_601;
wire sig_602;
wire sig_605;
wire sig_607;
wire sig_608;
wire sig_610;
wire sig_611;
wire sig_612;
wire sig_615;
wire sig_616;
wire sig_617;
wire sig_618;
wire sig_619;
wire sig_620;
wire sig_621;
wire sig_623;
wire sig_624;
wire sig_625;
wire sig_626;
wire sig_628;
wire sig_629;
wire sig_630;
wire sig_631;
wire sig_632;
wire sig_634;
wire sig_635;
wire sig_636;
wire sig_637;
wire sig_639;
wire sig_640;
wire sig_641;
wire sig_642;
wire sig_643;
wire sig_645;
wire sig_646;
wire sig_647;
wire sig_648;
wire sig_649;
wire sig_650;
wire sig_651;
wire sig_652;
wire sig_653;
wire sig_654;
wire sig_655;
wire sig_656;
wire sig_657;
wire sig_658;
wire sig_662;
wire sig_663;
wire sig_664;
wire sig_665;
wire sig_666;
wire sig_667;
wire sig_669;
wire sig_670;
wire sig_671;
wire sig_673;
wire sig_674;
wire sig_675;
wire sig_676;
wire sig_679;
wire sig_681;
wire sig_683;
wire sig_684;
wire sig_685;
wire sig_686;
wire sig_687;
wire sig_688;
wire sig_691;
wire sig_692;
wire sig_693;
wire sig_695;
wire sig_697;
wire sig_698;
wire sig_699;
wire sig_701;
wire sig_702;
wire sig_703;
wire sig_704;
wire sig_706;
wire sig_707;
wire sig_709;
wire sig_710;
wire sig_711;
wire sig_712;
wire sig_714;
wire sig_715;
wire sig_716;
wire sig_717;
wire sig_718;
wire sig_720;
wire sig_722;
wire sig_723;
wire sig_724;
wire sig_725;
wire sig_726;
wire sig_727;
wire sig_728;
wire sig_729;
wire sig_730;
wire sig_731;
wire sig_732;
wire sig_734;
wire sig_735;
wire sig_737;
wire sig_738;
wire sig_739;
wire sig_740;
wire sig_741;
wire sig_742;
wire sig_743;
wire sig_744;
wire sig_746;
wire sig_747;
wire sig_748;
wire sig_749;
wire sig_750;
wire sig_751;
wire sig_752;
wire sig_753;
wire sig_754;
wire sig_755;
wire sig_756;
wire sig_757;
wire sig_758;
wire sig_759;
wire sig_760;
wire sig_761;
wire sig_762;
wire sig_764;
wire sig_765;
wire sig_766;
wire sig_767;
wire sig_768;
wire sig_770;
wire sig_771;
wire sig_772;
wire sig_773;
wire sig_774;
wire sig_776;
wire sig_781;
wire sig_782;
wire sig_783;
wire sig_784;
wire sig_785;
wire sig_786;
wire sig_787;
wire sig_788;
wire sig_790;
wire sig_794;
wire sig_797;
wire sig_798;
wire sig_799;
wire sig_800;
wire sig_801;
wire sig_802;
wire sig_805;
wire sig_806;
wire sig_807;
wire sig_809;
wire sig_812;
wire sig_813;
wire sig_814;
wire sig_815;
wire sig_816;
wire sig_817;
wire sig_820;
wire sig_821;
wire sig_822;
wire sig_823;
wire sig_824;
wire sig_827;
wire sig_829;
wire sig_830;
wire sig_831;
wire sig_832;
wire sig_833;
wire sig_834;
wire sig_836;
wire sig_837;
wire sig_838;
wire sig_839;
wire sig_840;
wire sig_841;
wire sig_842;
wire sig_843;
wire sig_844;
wire sig_845;
wire sig_846;
wire sig_847;
wire sig_848;
wire sig_849;
wire sig_850;
wire sig_852;
wire sig_853;
wire sig_854;
wire sig_856;
wire sig_857;
wire sig_858;
wire sig_860;
wire sig_861;
wire sig_862;
wire sig_863;
wire sig_864;
wire sig_865;
wire sig_866;
wire sig_867;
wire sig_869;
wire sig_871;
wire sig_872;
wire sig_873;
wire sig_874;
wire sig_875;
wire sig_876;
wire sig_877;
wire sig_878;
wire sig_879;
wire sig_880;
wire sig_881;
wire sig_883;
wire sig_884;
wire sig_886;
wire sig_890;
wire sig_891;
wire sig_893;
wire sig_895;
wire sig_896;
wire sig_897;
wire sig_898;
wire sig_900;
wire sig_901;
wire sig_902;
wire sig_903;
wire sig_907;
wire sig_908;
wire sig_909;
wire sig_910;
wire sig_913;
wire sig_914;
wire sig_915;
wire sig_918;
wire sig_919;
wire sig_920;
wire sig_922;
wire sig_923;
wire sig_924;
wire sig_925;
wire sig_927;
wire sig_928;
wire sig_929;
wire sig_930;
wire sig_931;
wire sig_932;
wire sig_933;
wire sig_934;
wire sig_935;
wire sig_936;
wire sig_937;
wire sig_939;
wire sig_940;
wire sig_941;
wire sig_942;
wire sig_943;
wire sig_944;
wire sig_945;
wire sig_947;
wire sig_948;
wire sig_949;
wire sig_950;
wire sig_951;
wire sig_953;
wire sig_955;
wire sig_956;
wire sig_957;
wire sig_958;
wire sig_959;
wire sig_960;
wire sig_961;
wire sig_962;
wire sig_964;
wire sig_965;
wire sig_966;
wire sig_967;
wire sig_969;
wire sig_970;
wire sig_971;
wire sig_972;
wire sig_973;
wire sig_974;
wire sig_975;
wire sig_977;
wire sig_978;
wire sig_979;
wire sig_980;
wire sig_981;
wire sig_983;
wire sig_984;
wire sig_985;
wire sig_986;
wire sig_987;
wire sig_988;
wire sig_989;
wire sig_991;
wire sig_992;
wire sig_994;
wire sig_995;
wire sig_996;
wire sig_998;
wire sig_1000;
wire sig_1002;
wire sig_1004;
wire sig_1005;
wire sig_1006;
wire sig_1007;
wire sig_1009;
wire sig_1010;
wire sig_1011;
wire sig_1012;
wire sig_1013;
wire sig_1014;
wire sig_1015;
wire sig_1017;
wire sig_1018;
wire sig_1020;
wire sig_1021;
wire sig_1022;
wire sig_1023;
wire sig_1024;
wire sig_1025;
wire sig_1026;
wire sig_1027;
wire sig_1028;
wire sig_1029;
wire sig_1030;
wire sig_1032;
wire sig_1033;
wire sig_1034;
wire sig_1036;
wire sig_1037;
wire sig_1038;
wire sig_1039;
wire sig_1040;
wire sig_1041;
wire sig_1042;
wire sig_1045;
wire sig_1046;
wire sig_1047;
wire sig_1049;
wire sig_1050;
wire sig_1051;
wire sig_1053;
wire sig_1054;
wire sig_1055;
wire sig_1056;
wire sig_1058;
wire sig_1059;
wire sig_1060;
wire sig_1061;
wire sig_1062;
wire sig_1063;
wire sig_1065;
wire sig_1066;
wire sig_1068;
wire sig_1069;
wire sig_1070;
wire sig_1072;
wire sig_1073;
wire sig_1074;
wire sig_1076;
wire sig_1078;
wire sig_1079;
wire sig_1080;
wire sig_1082;
wire sig_1084;
wire sig_1085;
wire sig_1086;
wire sig_1087;
wire sig_1088;
wire sig_1089;
wire sig_1090;
wire sig_1091;
wire sig_1092;
wire sig_1093;
wire sig_1094;
wire sig_1095;
wire sig_1096;
wire sig_1098;
wire sig_1100;
wire sig_1102;
wire sig_1103;
wire sig_1105;
wire sig_1106;
wire sig_1107;
wire sig_1108;
wire sig_1109;
wire sig_1111;
wire sig_1112;
wire sig_1113;
wire sig_1114;
wire sig_1115;
wire sig_1117;
wire sig_1119;
wire sig_1120;
wire sig_1121;
wire sig_1122;
wire sig_1123;
wire sig_1124;
wire sig_1125;
wire sig_1126;
wire sig_1127;
wire sig_1129;
wire sig_1130;
wire sig_1131;
wire sig_1132;
wire sig_1133;
wire sig_1134;
wire sig_1135;
wire sig_1136;
wire sig_1137;
wire sig_1139;
wire sig_1140;
wire sig_1141;
wire sig_1142;
wire sig_1145;
wire sig_1146;
wire sig_1147;
wire sig_1148;
wire sig_1149;
wire sig_1150;
wire sig_1151;
wire sig_1152;
wire sig_1153;
wire sig_1154;
wire sig_1155;
wire sig_1156;
wire sig_1158;
wire sig_1159;
wire sig_1160;
wire sig_1161;
wire sig_1162;
wire sig_1163;
wire sig_1164;
wire sig_1165;
wire sig_1166;
wire sig_1167;
wire sig_1169;
wire sig_1170;
wire sig_1171;
wire sig_1172;
wire sig_1174;
wire sig_1175;
wire sig_1176;
wire sig_1177;
wire sig_1178;
wire sig_1180;
wire sig_1181;
wire sig_1182;
wire sig_1183;
wire sig_1185;
wire sig_1186;
wire sig_1187;
wire sig_1188;
wire sig_1189;
wire sig_1190;
wire sig_1191;
wire sig_1192;
wire sig_1193;
wire sig_1194;
wire sig_1195;
wire sig_1196;
wire sig_1197;
wire sig_1199;
wire sig_1200;
wire sig_1201;
wire sig_1202;
wire sig_1203;
wire sig_1204;
wire sig_1205;
wire sig_1206;
wire sig_1207;
wire sig_1209;
wire sig_1210;
wire sig_1213;
wire sig_1214;
wire sig_1215;
wire sig_1216;
wire sig_1218;
wire sig_1219;
wire sig_1220;
wire sig_1221;
wire sig_1222;
wire sig_1223;
wire sig_1225;
wire sig_1226;
wire sig_1227;
wire sig_1231;
wire sig_1232;
wire sig_1233;
wire sig_1234;
wire sig_1235;
wire sig_1237;
wire sig_1238;
wire sig_1240;
wire sig_1242;
wire sig_1244;
wire sig_1245;
wire sig_1246;
wire sig_1247;
wire sig_1248;
wire sig_1250;
wire sig_1251;
wire sig_1252;
wire sig_1253;
wire sig_1254;
wire sig_1256;
wire sig_1258;
wire sig_1259;
wire sig_1260;
wire sig_1262;
wire sig_1264;
wire sig_1266;
wire sig_1267;
wire sig_1268;
wire sig_1269;
wire sig_1270;
wire sig_1271;
wire sig_1272;
wire sig_1273;
wire sig_1274;
wire sig_1275;
wire sig_1277;
wire sig_1280;
wire sig_1281;
wire sig_1282;
wire sig_1283;
wire sig_1284;
wire sig_1285;
wire sig_1286;
wire sig_1287;
wire sig_1288;
wire sig_1289;
wire sig_1290;
wire sig_1291;
wire sig_1292;
wire sig_1293;
wire sig_1295;
wire sig_1296;
wire sig_1297;
wire sig_1299;
wire sig_1300;
wire sig_1301;
wire sig_1302;
wire sig_1303;
wire sig_1304;
wire sig_1305;
wire sig_1306;
wire sig_1307;
wire sig_1308;
wire sig_1309;
wire sig_1310;
wire sig_1311;
wire sig_1312;
wire sig_1313;
wire sig_1314;
wire sig_1316;
wire sig_1317;
wire sig_1318;
wire sig_1319;
wire sig_1320;
wire sig_1321;
wire sig_1323;
wire sig_1324;
wire sig_1325;
wire sig_1327;
wire sig_1328;
wire sig_1329;
wire sig_1330;
wire sig_1331;
wire sig_1332;
wire sig_1335;
wire sig_1337;
wire sig_1338;
wire sig_1339;
wire sig_1340;
wire sig_1342;
wire sig_1343;
wire sig_1344;
wire sig_1345;
wire sig_1346;
wire sig_1347;
wire sig_1349;
wire sig_1350;
wire sig_1351;
wire sig_1352;
wire sig_1353;
wire sig_1354;
wire sig_1355;
wire sig_1356;
wire sig_1357;
wire sig_1359;
wire sig_1360;
wire sig_1361;
wire sig_1362;
wire sig_1363;
wire sig_1364;
wire sig_1365;
wire sig_1366;
wire sig_1367;
wire sig_1368;
wire sig_1369;
wire sig_1370;
wire sig_1371;
wire sig_1372;
wire sig_1374;
wire sig_1377;
wire sig_1379;
wire sig_1380;
wire sig_1382;
wire sig_1383;
wire sig_1384;
wire sig_1385;
wire sig_1386;
wire sig_1387;
wire sig_1388;
wire sig_1389;
wire sig_1390;
wire sig_1391;
wire sig_1393;
wire sig_1394;
wire sig_1395;
wire sig_1397;
wire sig_1398;
wire sig_1400;
wire sig_1401;
wire sig_1402;
wire sig_1403;
wire sig_1404;
wire sig_1405;
wire sig_1406;
wire sig_1407;
wire sig_1408;
wire sig_1409;
wire sig_1410;
wire sig_1411;
wire sig_1412;
wire sig_1413;
wire sig_1414;
wire sig_1415;
wire sig_1416;
wire sig_1417;
wire sig_1419;
wire sig_1421;
wire sig_1422;
wire sig_1423;
wire sig_1424;
wire sig_1425;
wire sig_1427;
wire sig_1428;
wire sig_1429;
wire sig_1430;
wire sig_1431;
wire sig_1432;
wire sig_1433;
wire sig_1435;
wire sig_1436;
wire sig_1437;
wire sig_1438;
wire sig_1439;
wire sig_1440;
wire sig_1441;
wire sig_1442;
wire sig_1443;
wire sig_1444;
wire sig_1447;
wire sig_1449;
wire sig_1450;
wire sig_1451;
wire sig_1452;
wire sig_1454;
wire sig_1455;
wire sig_1456;
wire sig_1457;
wire sig_1458;
wire sig_1459;
wire sig_1461;
wire sig_1462;
wire sig_1464;
wire sig_1465;
wire sig_1467;
wire sig_1468;
wire sig_1469;
wire sig_1471;
wire sig_1472;
wire sig_1473;
wire sig_1474;
wire sig_1475;
wire sig_1477;
wire sig_1478;
wire sig_1479;
wire sig_1481;
wire sig_1483;
wire sig_1484;
wire sig_1485;
wire sig_1489;
wire sig_1490;
wire sig_1491;
wire sig_1492;
wire sig_1493;
wire sig_1497;
wire sig_1498;
wire sig_1499;
wire sig_1500;
wire sig_1501;
wire sig_1502;
wire sig_1503;
wire sig_1504;
wire sig_1505;
wire sig_1506;
wire sig_1507;
wire sig_1508;
wire sig_1509;
wire sig_1510;
wire sig_1511;
wire sig_1512;
wire sig_1513;
wire sig_1514;
wire sig_1515;
wire sig_1516;
wire sig_1517;
wire sig_1518;
wire sig_1519;
wire sig_1520;
wire sig_1521;
wire sig_1522;
wire sig_1523;
wire sig_1524;
wire sig_1525;
wire sig_1526;
wire sig_1527;
wire sig_1528;
wire sig_1529;
wire sig_1530;
wire sig_1531;
wire sig_1532;
wire sig_1533;
wire sig_1534;
wire sig_1535;
wire sig_1536;
wire sig_1537;
wire sig_1538;
wire sig_1539;
wire sig_1540;
wire sig_1541;
wire sig_1542;
wire sig_1543;
wire sig_1544;
wire sig_1545;
wire sig_1546;
wire sig_1547;
wire sig_1548;
wire sig_1549;
wire sig_1550;
wire sig_1551;
wire sig_1552;
wire sig_1553;
wire sig_1554;
wire sig_1555;
wire sig_1556;
wire sig_1557;
wire sig_1558;
wire sig_1559;
wire sig_1560;
wire sig_1561;
wire sig_1562;
wire sig_1563;
wire sig_1564;
wire sig_1565;

assign sig_32 = A[8] & B[6];
assign sig_33 = A[9] & B[5];
assign sig_34 = A[11] & B[14];
assign sig_36 = A[5] & B[15];
assign sig_37 = A[10] & B[3];
assign sig_38 = A[11] & B[11];
assign sig_39 = A[5] & B[9];
assign sig_40 = A[15] & B[13];
assign sig_41 = A[11] & B[0];
assign sig_42 = A[8] & B[8];
assign sig_43 = A[12] & B[13];
assign sig_44 = A[2] & B[12];
assign sig_45 = A[4] & B[11];
assign sig_46 = A[7] & B[6];
assign sig_47 = A[15] & B[8];
assign sig_49 = A[12] & B[1];
assign sig_50 = A[6] & B[15];
assign sig_52 = A[0] & A[4];
assign sig_54 = A[4] & B[9];
assign sig_55 = A[15] & B[14];
assign sig_56 = A[8] & B[11];
assign sig_57 = A[10] & B[14];
assign sig_58 = A[9] & B[4];
assign sig_59 = A[11] & B[7];
assign sig_60 = A[3] & B[11];
assign sig_62 = A[12] & B[11];
assign sig_64 = A[6] & B[13];
assign sig_66 = A[0] & B[13];
assign sig_67 = A[2] & B[15];
assign sig_69 = A[8] & B[0];
assign sig_70 = A[9] & B[8];
assign sig_71 = A[3] & B[12];
assign sig_72 = A[9] & B[13];
assign sig_73 = A[14] & B[10];
assign sig_74 = A[1] & B[10];
assign sig_75 = A[6] & B[6];
assign sig_76 = A[11] & B[5];
assign sig_77 = A[8] & B[4];
assign sig_78 = A[13] & B[14];
assign sig_79 = A[12] & B[7];
assign sig_80 = A[7] & B[15];
assign sig_84 = A[8] & B[3];
assign sig_85 = A[3] & B[9];
assign sig_86 = A[4] & B[14];
assign sig_87 = A[6] & B[8];
assign sig_88 = A[10] & B[13];
assign sig_90 = A[13] & B[0];
assign sig_91 = A[6] & B[11];
assign sig_92 = A[5] & B[6];
assign sig_93 = A[15] & B[7];
assign sig_94 = A[12] & B[5];
assign sig_95 = A[14] & B[6];
assign sig_96 = A[1] & B[15];
assign sig_97 = A[11] & B[12];
assign sig_98 = A[8] & B[15];
assign sig_99 = A[3] & B[15];
assign sig_100 = A[2] & B[10];
assign sig_101 = A[2] & B[9];
assign sig_102 = A[5] & B[14];
assign sig_103 = A[11] & B[4];
assign sig_104 = A[11] & B[1];
assign sig_105 = A[12] & B[14];
assign sig_107 = A[15] & B[6];
assign sig_108 = A[10] & B[12];
assign sig_109 = A[7] & B[8];
assign sig_110 = A[1] & B[12];
assign sig_111 = A[12] & B[0];
assign sig_112 = A[3] & B[10];
assign sig_115 = A[11] & B[2];
assign sig_117 = A[10] & B[4];
assign sig_119 = A[7] & B[14];
assign sig_120 = A[9] & B[15];
assign sig_123 = A[1] & B[9];
assign sig_124 = sig_101 & sig_74;
assign sig_125 = A[0] & B[14];
assign sig_126 = A[0] & B[11];
assign sig_127 = A[10] & B[2];
assign sig_128 = A[12] & B[9];
assign sig_129 = A[6] & B[5];
assign sig_131 = A[8] & B[13];
assign sig_132 = A[10] & B[8];
assign sig_133 = A[9] & B[12];
assign sig_134 = A[10] & B[15];
assign sig_137 = A[4] & B[10];
assign sig_138 = A[13] & B[4];
assign sig_140 = A[6] & B[14];
assign sig_141 = A[1] & B[14];
assign sig_142 = A[5] & B[7];
assign sig_143 = sig_97 & sig_88;
assign sig_145 = A[8] & B[12];
assign sig_146 = A[4] & B[13];
assign sig_147 = A[10] & B[5];
assign sig_148 = A[11] & B[8];
assign sig_149 = sig_85 & sig_100;
assign sig_150 = A[5] & B[10];
assign sig_151 = A[9] & B[2];
assign sig_152 = A[7] & B[5];
assign sig_153 = sig_88 ^ sig_105;
assign sig_154 = A[12] & B[4];
assign sig_155 = A[5] & B[13];
assign sig_157 = A[13] & B[10];
assign sig_158 = A[9] & B[14];
assign sig_160 = sig_75 ^ sig_142;
assign sig_161 = A[11] & B[15];
assign sig_162 = A[6] & B[7];
assign sig_163 = sig_108 & sig_72;
assign sig_164 = A[15] & B[11];
assign sig_168 = A[14] & B[4];
assign sig_169 = A[2] & B[11];
assign sig_170 = sig_54 & sig_112;
assign sig_171 = A[2] & B[14];
assign sig_173 = A[8] & B[2];
assign sig_174 = A[8] & B[5];
assign sig_176 = A[15] & B[12];
assign sig_177 = A[3] & B[13];
assign sig_179 = A[15] & B[9];
assign sig_180 = A[12] & B[15];
assign sig_181 = sig_46 ^ sig_162;
assign sig_182 = A[6] & B[10];
assign sig_183 = A[15] & B[10];
assign sig_186 = A[8] & B[14];
assign sig_187 = A[5] & B[11];
assign sig_188 = A[3] & B[14];
assign sig_189 = A[10] & B[1];
assign sig_191 = sig_133 & sig_131;
assign sig_194 = A[14] & B[12];
assign sig_195 = A[1] & B[11];
assign sig_196 = A[15] & B[3];
assign sig_197 = sig_90 ^ sig_49;
assign sig_198 = A[7] & B[10];
assign sig_201 = A[2] & B[13];
assign sig_203 = sig_101 ^ sig_74;
assign sig_206 = A[13] & B[15];
assign sig_208 = A[4] & B[7];
assign sig_210 = sig_111 ^ sig_104;
assign sig_211 = A[13] & B[11];
assign sig_212 = A[14] & B[2];
assign sig_213 = A[1] & B[13];
assign sig_214 = A[15] & B[2];
assign sig_215 = A[13] & B[12];
assign sig_217 = sig_46 & sig_162;
assign sig_218 = A[14] & B[15];
assign sig_219 = A[8] & B[10];
assign sig_220 = sig_133 ^ sig_131;
assign sig_223 = A[10] & B[9];
assign sig_224 = A[14] & B[11];
assign sig_225 = A[15] & B[5];
assign sig_226 = A[9] & B[7];
assign sig_229 = A[12] & B[12];
assign sig_230 = A[13] & B[3];
assign sig_233 = A[9] & B[10];
assign sig_234 = sig_37 ^ sig_58;
assign sig_235 = A[13] & B[2];
assign sig_236 = sig_54 ^ sig_112;
assign sig_239 = sig_75 & sig_142;
assign sig_240 = A[10] & B[7];
assign sig_244 = sig_108 ^ sig_72;
assign sig_245 = A[14] & B[3];
assign sig_246 = A[9] & B[9];
assign sig_247 = A[13] & B[1];
assign sig_248 = A[14] & B[7];
assign sig_249 = A[15] & B[0];
assign sig_250 = A[11] & B[10];
assign sig_252 = A[12] & B[2];
assign sig_253 = A[6] & B[12];
assign sig_254 = A[13] & B[6];
assign sig_256 = A[4] & B[8];
assign sig_257 = sig_223 & sig_233;
assign sig_259 = A[11] & B[6];
assign sig_260 = sig_259 ^ sig_240;
assign sig_261 = sig_92 & sig_208;
assign sig_263 = sig_41 & sig_189;
assign sig_264 = sig_97 ^ sig_88;
assign sig_266 = sig_37 & sig_58;
assign sig_269 = sig_85 ^ sig_100;
assign sig_270 = A[8] & B[9];
assign sig_271 = A[14] & B[1];
assign sig_272 = A[13] & B[7];
assign sig_273 = sig_215 & sig_43;
assign sig_274 = A[14] & B[14];
assign sig_276 = A[7] & B[7];
assign sig_278 = A[13] & B[9];
assign sig_279 = A[5] & B[8];
assign sig_281 = A[11] & B[3];
assign sig_283 = A[13] & B[5];
assign sig_284 = A[15] & B[15];
assign sig_285 = A[4] & B[15];
assign sig_286 = A[14] & B[0];
assign sig_287 = A[10] & B[10];
assign sig_288 = A[13] & B[13];
assign sig_290 = A[7] & B[12];
assign sig_291 = A[14] & B[8];
assign sig_292 = A[12] & B[6];
assign sig_295 = A[0] & B[12];
assign sig_297 = A[10] & B[6];
assign sig_299 = sig_292 ^ sig_59;
assign sig_300 = A[7] & B[13];
assign sig_301 = A[8] & B[7];
assign sig_302 = A[15] & B[1];
assign sig_303 = A[12] & B[3];
assign sig_304 = A[9] & B[11];
assign sig_305 = sig_71 & sig_148;
assign sig_306 = A[7] & B[9];
assign sig_308 = A[14] & B[13];
assign sig_309 = A[13] & B[8];
assign sig_311 = A[4] & B[12];
assign sig_312 = A[14] & B[9];
assign sig_315 = A[9] & B[6];
assign sig_316 = sig_254 ^ sig_79;
assign sig_317 = sig_119 & sig_220;
assign sig_318 = A[14] & B[5];
assign sig_319 = sig_90 & sig_49;
assign sig_320 = sig_132 & sig_299;
assign sig_321 = sig_215 ^ sig_43;
assign sig_324 = sig_39 ^ sig_137;
assign sig_326 = A[6] & B[9];
assign sig_328 = A[15] & B[4];
assign sig_329 = A[7] & B[4];
assign sig_330 = A[11] & B[9];
assign sig_331 = sig_39 & sig_137;
assign sig_332 = A[7] & B[11];
assign sig_333 = A[9] & B[3];
assign sig_334 = sig_249 ^ sig_271;
assign sig_335 = A[10] & B[11];
assign sig_336 = sig_111 & sig_104;
assign sig_337 = A[0] & B[15];
assign sig_338 = sig_107 ^ sig_248;
assign sig_339 = A[3] & B[8];
assign sig_340 = A[11] & B[13];
assign sig_341 = A[12] & B[8];
assign sig_343 = sig_291 & sig_93;
assign sig_345 = A[12] & B[10];
assign sig_346 = A[5] & B[12];
assign sig_347 = sig_260 ^ sig_70;
assign sig_348 = sig_84 & sig_329;
assign sig_349 = sig_270 ^ sig_198;
assign sig_351 = sig_174 & sig_234;
assign sig_352 = sig_148 & sig_316;
assign sig_353 = sig_194 ^ sig_288;
assign sig_354 = sig_110 & sig_66;
assign sig_355 = sig_286 ^ sig_247;
assign sig_356 = sig_333 ^ sig_77;
assign sig_359 = sig_326 & sig_150;
assign sig_360 = sig_249 & sig_271;
assign sig_361 = sig_95 ^ sig_272;
assign sig_364 = sig_176 ^ sig_308;
assign sig_365 = sig_253 & sig_155;
assign sig_366 = sig_93 ^ sig_291;
assign sig_367 = sig_306 ^ sig_182;
assign sig_368 = sig_311 & sig_177;
assign sig_369 = sig_328 ^ sig_318;
assign sig_371 = sig_324 ^ sig_60;
assign sig_372 = sig_152 & sig_356;
assign sig_373 = sig_306 & sig_182;
assign sig_374 = sig_91 & sig_349;
assign sig_375 = sig_286 & sig_247;
assign sig_376 = sig_110 ^ sig_66;
assign sig_378 = sig_197 ^ sig_115;
assign sig_379 = sig_223 ^ sig_233;
assign sig_380 = sig_330 ^ sig_287;
assign sig_381 = sig_349 ^ sig_91;
assign sig_382 = sig_290 & sig_64;
assign sig_383 = sig_40 ^ sig_274;
assign sig_384 = sig_346 & sig_146;
assign sig_385 = sig_270 & sig_198;
assign sig_388 = sig_220 ^ sig_119;
assign sig_390 = sig_123 & sig_52;
assign sig_391 = sig_254 & sig_79;
assign sig_393 = sig_246 ^ sig_219;
assign sig_394 = sig_128 ^ sig_250;
assign sig_395 = sig_364 ^ sig_78;
assign sig_396 = sig_44 & sig_213;
assign sig_397 = sig_367 ^ sig_187;
assign sig_398 = sig_318 & sig_328;
assign sig_401 = sig_84 ^ sig_329;
assign sig_402 = sig_126 & sig_203;
assign sig_403 = sig_127 & sig_210;
assign sig_404 = sig_338 ^ sig_309;
assign sig_405 = sig_191 | sig_317;
assign sig_406 = sig_41 ^ sig_189;
assign sig_407 = sig_181 ^ sig_279;
assign sig_408 = sig_196 ^ sig_168;
assign sig_410 = sig_278 ^ sig_345;
assign sig_413 = sig_203 | sig_126;
assign sig_414 = sig_124 | sig_402;
assign sig_415 = sig_292 & sig_59;
assign sig_417 = sig_196 & sig_168;
assign sig_419 = sig_195 & sig_269;
assign sig_420 = sig_115 & sig_197;
assign sig_421 = sig_71 & sig_201;
assign sig_422 = sig_71 ^ sig_201;
assign sig_423 = sig_160 ^ sig_256;
assign sig_426 = sig_212 & sig_302;
assign sig_427 = sig_264 ^ sig_158;
assign sig_428 = sig_256 & sig_160;
assign sig_429 = sig_92 ^ sig_208;
assign sig_430 = sig_259 & sig_240;
assign sig_432 = sig_312 ^ sig_157;
assign sig_433 = sig_44 ^ sig_213;
assign sig_434 = sig_149 | sig_419;
assign sig_437 = sig_245 ^ sig_138;
assign sig_438 = sig_169 & sig_236;
assign sig_439 = sig_183 ^ sig_224;
assign sig_440 = sig_244 ^ sig_186;
assign sig_442 = sig_429 ^ sig_339;
assign sig_443 = sig_105 & sig_353;
assign sig_444 = sig_179 ^ sig_73;
assign sig_446 = sig_236 ^ sig_169;
assign sig_447 = sig_170 | sig_438;
assign sig_448 = sig_279 & sig_181;
assign sig_449 = sig_297 & sig_226;
assign sig_451 = sig_230 ^ sig_154;
assign sig_453 = sig_356 ^ sig_152;
assign sig_454 = sig_346 ^ sig_146;
assign sig_458 = sig_299 ^ sig_132;
assign sig_460 = sig_210 ^ sig_127;
assign sig_461 = sig_321 ^ sig_34;
assign sig_462 = sig_179 & sig_73;
assign sig_463 = sig_334 ^ sig_235;
assign sig_466 = sig_69 ^ sig_305;
assign sig_467 = sig_315 & sig_301;
assign sig_468 = sig_78 & sig_364;
assign sig_469 = sig_234 ^ sig_174;
assign sig_470 = sig_311 ^ sig_177;
assign sig_472 = sig_95 & sig_272;
assign sig_473 = sig_309 & sig_338;
assign sig_474 = sig_269 ^ sig_195;
assign sig_475 = sig_37 & sig_390;
assign sig_476 = sig_230 & sig_154;
assign sig_477 = sig_283 & sig_408;
assign sig_481 = sig_303 ^ sig_103;
assign sig_482 = sig_355 ^ sig_252;
assign sig_485 = sig_319 | sig_420;
assign sig_486 = sig_341 & sig_361;
assign sig_487 = sig_245 & sig_138;
assign sig_488 = sig_47 ^ sig_343;
assign sig_489 = sig_32 & sig_276;
assign sig_490 = sig_339 & sig_429;
assign sig_491 = sig_32 ^ sig_276;
assign sig_492 = sig_147 & sig_481;
assign sig_493 = sig_145 & sig_300;
assign sig_494 = sig_380 ^ sig_304;
assign sig_495 = sig_281 ^ sig_117;
assign sig_496 = sig_290 ^ sig_64;
assign sig_497 = sig_107 & sig_248;
assign sig_498 = sig_335 & sig_394;
assign sig_500 = sig_332 & sig_393;
assign sig_501 = sig_336 | sig_403;
assign sig_502 = sig_224 & sig_183;
assign sig_503 = sig_315 ^ sig_301;
assign sig_504 = sig_34 & sig_321;
assign sig_505 = sig_145 ^ sig_300;
assign sig_506 = sig_253 ^ sig_155;
assign sig_507 = sig_401 | sig_129;
assign sig_508 = sig_281 & sig_117;
assign sig_509 = sig_266 | sig_351;
assign sig_510 = sig_304 & sig_380;
assign sig_511 = sig_56 & sig_379;
assign sig_512 = sig_33 & sig_495;
assign sig_513 = sig_176 & sig_308;
assign sig_514 = sig_394 ^ sig_335;
assign sig_515 = sig_513 | sig_468;
assign sig_516 = sig_302 ^ sig_212;
assign sig_517 = sig_128 & sig_250;
assign sig_518 = sig_353 ^ sig_105;
assign sig_519 = sig_246 & sig_219;
assign sig_520 = sig_186 & sig_244;
assign sig_521 = sig_303 & sig_103;
assign sig_522 = B[7] | sig_442;
assign sig_523 = sig_297 ^ sig_226;
assign sig_524 = sig_70 & sig_260;
assign sig_525 = sig_343 & sig_47;
assign sig_526 = sig_94 & sig_437;
assign sig_527 = sig_194 & sig_288;
assign sig_529 = sig_379 ^ sig_56;
assign sig_530 = sig_451 ^ sig_76;
assign sig_532 = sig_62 & sig_432;
assign sig_533 = sig_410 ^ sig_38;
assign sig_534 = sig_274 & sig_40;
assign sig_535 = sig_330 & sig_287;
assign sig_536 = sig_87 & sig_491;
assign sig_537 = sig_158 & sig_264;
assign sig_538 = sig_214 ^ sig_426;
assign sig_539 = sig_446 & sig_434;
assign sig_540 = sig_164 & sig_502;
assign sig_541 = sig_393 ^ sig_332;
assign sig_542 = sig_437 ^ sig_94;
assign sig_544 = sig_519 | sig_500;
assign sig_545 = sig_432 ^ sig_62;
assign sig_546 = sig_76 & sig_451;
assign sig_548 = sig_474 ^ sig_414;
assign sig_549 = sig_333 & sig_77;
assign sig_550 = sig_38 & sig_410;
assign sig_551 = sig_391 | sig_352;
assign sig_552 = sig_295 & sig_548;
assign sig_553 = sig_252 & sig_355;
assign sig_554 = sig_140 & sig_505;
assign sig_555 = sig_69 & B[6];
assign sig_556 = sig_474 & sig_414;
assign sig_557 = sig_312 & sig_157;
assign sig_558 = sig_316 ^ sig_148;
assign sig_559 = sig_257 | sig_511;
assign sig_560 = sig_476 | sig_546;
assign sig_561 = sig_326 ^ sig_150;
assign sig_563 = sig_109 & sig_503;
assign sig_564 = sig_229 & sig_340;
assign sig_565 = sig_129 & sig_401;
assign sig_567 = sig_446 ^ sig_434;
assign sig_568 = sig_229 ^ sig_340;
assign sig_570 = sig_495 ^ sig_33;
assign sig_571 = sig_415 | sig_320;
assign sig_572 = sig_235 & sig_334;
assign sig_573 = sig_60 & sig_324;
assign sig_574 = sig_278 & sig_345;
assign sig_577 = sig_517 | sig_498;
assign sig_578 = sig_361 ^ sig_341;
assign sig_579 = sig_413 | sig_390;
assign sig_580 = sig_494 & sig_559;
assign sig_581 = sig_331 | sig_573;
assign sig_582 = sig_481 ^ sig_147;
assign sig_585 = sig_487 | sig_526;
assign sig_586 = sig_538 ^ sig_542;
assign sig_587 = sig_522 ^ sig_428;
assign sig_588 = sig_45 & sig_561;
assign sig_589 = sig_398 & sig_578;
assign sig_590 = sig_371 ^ sig_447;
assign sig_592 = sig_430 | sig_524;
assign sig_594 = sig_508 ^ sig_512;
assign sig_595 = sig_535 | sig_510;
assign sig_596 = sig_188 & sig_454;
assign sig_597 = sig_433 ^ sig_125;
assign sig_598 = sig_561 ^ sig_45;
assign sig_599 = sig_598 ^ sig_581;
assign sig_601 = sig_514 & sig_595;
assign sig_602 = sig_359 | sig_588;
assign sig_605 = sig_408 ^ sig_283;
assign sig_607 = sig_187 & sig_367;
assign sig_608 = sig_523 ^ sig_42;
assign sig_610 = sig_171 & sig_470;
assign sig_611 = sig_557 | sig_532;
assign sig_612 = sig_422 ^ sig_141;
assign sig_615 = sig_560 ^ sig_347;
assign sig_616 = sig_533 & sig_577;
assign sig_617 = sig_373 | sig_607;
assign sig_618 = sig_529 & sig_544;
assign sig_619 = sig_397 ^ sig_602;
assign sig_620 = sig_521 | sig_492;
assign sig_621 = sig_585 ^ sig_458;
assign sig_623 = sig_467 | sig_563;
assign sig_624 = sig_514 ^ sig_595;
assign sig_625 = sig_173 & sig_466;
assign sig_626 = sig_560 & sig_347;
assign sig_628 = sig_620 ^ sig_608;
assign sig_629 = sig_472 | sig_486;
assign sig_630 = sig_503 ^ sig_109;
assign sig_631 = sig_574 | sig_550;
assign sig_632 = sig_141 & sig_422;
assign sig_634 = sig_360 | sig_572;
assign sig_635 = sig_470 ^ sig_171;
assign sig_636 = sig_556 | sig_552;
assign sig_637 = sig_417 | sig_477;
assign sig_639 = sig_381 ^ sig_617;
assign sig_640 = sig_545 & sig_631;
assign sig_641 = sig_506 ^ sig_86;
assign sig_642 = sig_385 | sig_374;
assign sig_643 = sig_529 ^ sig_544;
assign sig_645 = sig_612 & sig_599;
assign sig_646 = sig_421 | sig_632;
assign sig_647 = sig_494 ^ sig_559;
assign sig_648 = sig_151 & sig_406;
assign sig_649 = sig_49 & sig_155;
assign sig_650 = sig_482 & sig_485;
assign sig_651 = sig_491 ^ sig_87;
assign sig_652 = sig_497 | sig_473;
assign sig_653 = sig_489 | sig_536;
assign sig_654 = sig_125 & sig_433;
assign sig_655 = sig_454 ^ sig_188;
assign sig_656 = sig_493 | sig_554;
assign sig_657 = sig_406 ^ sig_151;
assign sig_658 = sig_496 ^ sig_102;
assign sig_662 = sig_217 | sig_448;
assign sig_663 = sig_375 | sig_553;
assign sig_664 = sig_218 & sig_534;
assign sig_665 = sig_597 & sig_590;
assign sig_666 = sig_396 | sig_654;
assign sig_667 = sig_545 ^ sig_631;
assign sig_669 = sig_522 & sig_442;
assign sig_670 = sig_505 ^ sig_140;
assign sig_671 = sig_509 ^ sig_651;
assign sig_673 = sig_534 ^ sig_218;
assign sig_674 = sig_214 & sig_426;
assign sig_675 = sig_594 ^ sig_630;
assign sig_676 = sig_621 ^ sig_592;
assign sig_679 = sig_102 & sig_496;
assign sig_681 = sig_548 ^ sig_295;
assign sig_683 = sig_444 ^ sig_211;
assign sig_684 = sig_384 | sig_596;
assign sig_685 = sig_533 ^ sig_577;
assign sig_686 = sig_516 & sig_634;
assign sig_687 = sig_382 | sig_679;
assign sig_688 = sig_239 | sig_428;
assign sig_691 = sig_163 | sig_520;
assign sig_692 = sig_598 & sig_581;
assign sig_693 = sig_86 & sig_506;
assign sig_695 = sig_567 ^ sig_376;
assign sig_697 = sig_261 | sig_490;
assign sig_698 = sig_211 & sig_444;
assign sig_699 = sig_368 | sig_610;
assign sig_701 = sig_143 | sig_537;
assign sig_702 = sig_365 | sig_693;
assign sig_703 = sig_371 & sig_447;
assign sig_704 = sig_263 | sig_648;
assign sig_706 = sig_683 ^ sig_611;
assign sig_707 = sig_349 & sig_299;
assign sig_709 = sig_398 ^ sig_578;
assign sig_710 = sig_407 & sig_684;
assign sig_711 = sig_555 | sig_625;
assign sig_712 = sig_542 & sig_538;
assign sig_714 = sig_366 ^ sig_652;
assign sig_715 = sig_381 & sig_617;
assign sig_716 = sig_378 ^ sig_501;
assign sig_717 = sig_667 ^ sig_427;
assign sig_718 = sig_55 ^ sig_673;
assign sig_720 = sig_568 ^ sig_57;
assign sig_722 = sig_273 | sig_504;
assign sig_723 = sig_378 & sig_501;
assign sig_724 = sig_57 & sig_568;
assign sig_725 = sig_482 ^ sig_485;
assign sig_726 = sig_397 & sig_602;
assign sig_727 = sig_619 ^ sig_635;
assign sig_728 = sig_549 | sig_372;
assign sig_729 = sig_440 & sig_685;
assign sig_730 = sig_164 ^ sig_502;
assign sig_731 = sig_685 ^ sig_440;
assign sig_732 = sig_460 & sig_704;
assign sig_734 = sig_616 | sig_729;
assign sig_735 = sig_527 | sig_443;
assign sig_737 = sig_42 & sig_523;
assign sig_738 = sig_652 & sig_366;
assign sig_739 = sig_463 ^ sig_663;
assign sig_740 = sig_653 & sig_675;
assign sig_741 = sig_683 & sig_611;
assign sig_742 = sig_624 ^ sig_388;
assign sig_743 = sig_639 ^ sig_655;
assign sig_744 = sig_551 & sig_709;
assign sig_746 = sig_516 ^ sig_634;
assign sig_747 = sig_590 ^ sig_597;
assign sig_748 = sig_462 | sig_698;
assign sig_749 = sig_404 ^ sig_629;
assign sig_750 = sig_720 & sig_706;
assign sig_751 = sig_662 & sig_671;
assign sig_752 = sig_439 & sig_748;
assign sig_753 = sig_658 & sig_643;
assign sig_754 = sig_647 ^ sig_670;
assign sig_755 = sig_376 & sig_567;
assign sig_756 = sig_585 & sig_458;
assign sig_757 = sig_587 | sig_153;
assign sig_758 = sig_741 | sig_750;
assign sig_759 = sig_673 & sig_55;
assign sig_760 = sig_589 | sig_744;
assign sig_761 = sig_599 ^ sig_612;
assign sig_762 = sig_637 & sig_558;
assign sig_764 = sig_628 ^ sig_623;
assign sig_765 = sig_348 | sig_565;
assign sig_766 = sig_629 & sig_404;
assign sig_767 = sig_592 & sig_621;
assign sig_768 = sig_284 ^ sig_759;
assign sig_770 = sig_623 & sig_628;
assign sig_771 = sig_509 & sig_651;
assign sig_772 = sig_670 & sig_647;
assign sig_773 = sig_427 & sig_667;
assign sig_774 = sig_768 ^ sig_664;
assign sig_776 = sig_388 & sig_624;
assign sig_781 = sig_594 & sig_630;
assign sig_782 = sig_674 | sig_712;
assign sig_783 = sig_709 ^ sig_551;
assign sig_784 = sig_558 & sig_415;
assign sig_785 = sig_671 ^ sig_662;
assign sig_786 = sig_449 | sig_737;
assign sig_787 = sig_620 & sig_608;
assign sig_788 = sig_655 & sig_639;
assign sig_790 = sig_746 ^ sig_530;
assign sig_794 = sig_675 ^ sig_653;
assign sig_797 = sig_637 ^ sig_558;
assign sig_798 = sig_539 | sig_755;
assign sig_799 = sig_766 ^ sig_731;
assign sig_800 = sig_781 | sig_740;
assign sig_801 = sig_643 ^ sig_658;
assign sig_802 = sig_739 ^ sig_582;
assign sig_805 = sig_541 ^ sig_642;
assign sig_806 = sig_783 & sig_225;
assign sig_807 = sig_635 & sig_619;
assign sig_809 = sig_463 & sig_663;
assign sig_812 = sig_541 & sig_642;
assign sig_813 = sig_771 | sig_751;
assign sig_814 = sig_800 ^ sig_727;
assign sig_815 = sig_738 & sig_717;
assign sig_816 = sig_738 ^ sig_717;
assign sig_817 = sig_725 ^ sig_570;
assign sig_820 = sig_813 ^ sig_761;
assign sig_821 = sig_692 | sig_645;
assign sig_822 = sig_469 & sig_716;
assign sig_823 = sig_716 ^ sig_469;
assign sig_824 = sig_766 & sig_731;
assign sig_827 = sig_723 | sig_822;
assign sig_829 = sig_703 | sig_665;
assign sig_830 = sig_760 & sig_742;
assign sig_831 = sig_734 & sig_816;
assign sig_832 = sig_760 ^ sig_742;
assign sig_833 = sig_765 & sig_423;
assign sig_834 = sig_730 ^ sig_518;
assign sig_836 = sig_797 ^ sig_571;
assign sig_837 = sig_605 ^ sig_782;
assign sig_838 = sig_715 | sig_788;
assign sig_839 = sig_817 & sig_827;
assign sig_840 = sig_728 ^ sig_407;
assign sig_841 = sig_674 & sig_233;
assign sig_842 = sig_676 & sig_837;
assign sig_843 = sig_657 ^ sig_711;
assign sig_844 = sig_710 & sig_587;
assign sig_845 = sig_728 & sig_407;
assign sig_846 = sig_439 ^ sig_748;
assign sig_847 = sig_530 & sig_746;
assign sig_848 = sig_765 ^ sig_423;
assign sig_849 = sig_657 & sig_711;
assign sig_850 = sig_460 ^ sig_704;
assign sig_852 = sig_726 | sig_807;
assign sig_853 = sig_756 | sig_767;
assign sig_854 = sig_800 & sig_727;
assign sig_856 = sig_706 ^ sig_720;
assign sig_857 = sig_821 & sig_814;
assign sig_858 = sig_518 & sig_730;
assign sig_860 = sig_618 | sig_753;
assign sig_861 = sig_580 | sig_772;
assign sig_862 = sig_564 | sig_724;
assign sig_863 = sig_605 & sig_782;
assign sig_864 = sig_664 & sig_768;
assign sig_865 = sig_688 & sig_840;
assign sig_866 = sig_525 ^ sig_856;
assign sig_867 = sig_641 & sig_805;
assign sig_869 = sig_570 & sig_725;
assign sig_871 = sig_848 ^ sig_697;
assign sig_872 = sig_812 | sig_867;
assign sig_873 = sig_601 | sig_776;
assign sig_874 = sig_697 & sig_848;
assign sig_875 = sig_284 & sig_759;
assign sig_876 = sig_840 ^ sig_688;
assign sig_877 = sig_817 ^ sig_827;
assign sig_878 = sig_832 ^ sig_861;
assign sig_879 = sig_582 & sig_739;
assign sig_880 = sig_225 ^ sig_783;
assign sig_881 = sig_813 & sig_761;
assign sig_883 = sig_845 | sig_865;
assign sig_884 = sig_815 | sig_831;
assign sig_886 = sig_461 & sig_846;
assign sig_890 = sig_875 | sig_864;
assign sig_891 = sig_640 | sig_773;
assign sig_893 = sig_836 & sig_369;
assign sig_895 = sig_786 & sig_615;
assign sig_896 = sig_853 & sig_801;
assign sig_897 = sig_891 & sig_866;
assign sig_898 = sig_669 | sig_844;
assign sig_900 = sig_571 & sig_797;
assign sig_901 = sig_820 ^ sig_829;
assign sig_902 = sig_752 | sig_886;
assign sig_903 = sig_854 | sig_857;
assign sig_907 = sig_814 ^ sig_821;
assign sig_908 = sig_707 & sig_339;
assign sig_909 = sig_615 ^ sig_786;
assign sig_910 = sig_540 | sig_858;
assign sig_913 = sig_853 ^ sig_801;
assign sig_914 = sig_686 | sig_847;
assign sig_915 = sig_626 | sig_895;
assign sig_918 = sig_913 ^ sig_872;
assign sig_919 = sig_880 & sig_893;
assign sig_920 = sig_799 ^ sig_873;
assign sig_922 = sig_787 | sig_770;
assign sig_923 = sig_805 ^ sig_641;
assign sig_924 = sig_861 & sig_832;
assign sig_925 = sig_915 ^ sig_923;
assign sig_927 = sig_714 ^ sig_920;
assign sig_928 = sig_749 & sig_806;
assign sig_929 = sig_707 & sig_908;
assign sig_930 = sig_922 ^ sig_743;
assign sig_931 = sig_650 | sig_869;
assign sig_932 = sig_816 ^ sig_734;
assign sig_933 = sig_525 & sig_856;
assign sig_934 = sig_488 ^ sig_932;
assign sig_935 = sig_872 & sig_913;
assign sig_936 = sig_749 ^ sig_806;
assign sig_937 = sig_453 & sig_850;
assign sig_939 = sig_809 | sig_879;
assign sig_940 = sig_838 & sig_925;
assign sig_941 = sig_898 & sig_681;
assign sig_942 = sig_880 ^ sig_893;
assign sig_943 = sig_884 ^ sig_701;
assign sig_944 = sig_749 & sig_724;
assign sig_945 = sig_896 | sig_935;
assign sig_947 = sig_732 | sig_937;
assign sig_948 = sig_873 & sig_799;
assign sig_949 = sig_863 | sig_842;
assign sig_950 = sig_369 ^ sig_836;
assign sig_951 = sig_829 & sig_820;
assign sig_953 = sig_843 ^ sig_507;
assign sig_955 = sig_883 ^ sig_747;
assign sig_956 = sig_837 ^ sig_676;
assign sig_957 = sig_802 & sig_931;
assign sig_958 = sig_866 ^ sig_891;
assign sig_959 = sig_850 ^ sig_453;
assign sig_960 = sig_798 & sig_955;
assign sig_961 = sig_902 & sig_834;
assign sig_962 = sig_833 | sig_874;
assign sig_964 = sig_507 & sig_843;
assign sig_965 = sig_395 ^ sig_910;
assign sig_966 = sig_962 ^ sig_695;
assign sig_967 = sig_762 | sig_900;
assign sig_969 = sig_846 ^ sig_461;
assign sig_970 = sig_852 & sig_930;
assign sig_971 = sig_967 & sig_754;
assign sig_972 = sig_910 & sig_395;
assign sig_973 = sig_884 & sig_701;
assign sig_974 = sig_950 & sig_949;
assign sig_975 = sig_849 | sig_964;
assign sig_977 = sig_898 ^ sig_681;
assign sig_978 = sig_586 & sig_914;
assign sig_979 = sig_877 ^ sig_785;
assign sig_980 = sig_955 ^ sig_798;
assign sig_981 = sig_834 ^ sig_902;
assign sig_983 = sig_933 | sig_897;
assign sig_984 = sig_707 ^ sig_908;
assign sig_985 = sig_790 ^ sig_939;
assign sig_986 = sig_120 & sig_943;
assign sig_987 = sig_790 & sig_939;
assign sig_988 = sig_903 ^ sig_699;
assign sig_989 = sig_922 & sig_743;
assign sig_991 = sig_785 & sig_877;
assign sig_992 = sig_758 & sig_969;
assign sig_994 = sig_846 & sig_475;
assign sig_995 = sig_977 ^ sig_579;
assign sig_996 = sig_586 ^ sig_914;
assign sig_998 = sig_883 & sig_747;
assign sig_1000 = sig_824 | sig_948;
assign sig_1002 = sig_636 & sig_966;
assign sig_1004 = sig_764 & sig_985;
assign sig_1005 = sig_945 & sig_687;
assign sig_1006 = sig_1000 ^ sig_691;
assign sig_1007 = sig_802 ^ sig_931;
assign sig_1009 = sig_909 & sig_996;
assign sig_1010 = sig_973 | sig_986;
assign sig_1011 = sig_915 & sig_923;
assign sig_1012 = sig_579 & sig_977;
assign sig_1013 = sig_878 & sig_936;
assign sig_1014 = sig_959 ^ sig_975;
assign sig_1015 = sig_944 & sig_153;
assign sig_1017 = sig_930 ^ sig_852;
assign sig_1018 = A[1] & sig_984;
assign sig_1020 = sig_830 | sig_924;
assign sig_1021 = sig_903 & sig_699;
assign sig_1022 = sig_932 & sig_488;
assign sig_1023 = sig_98 & sig_1006;
assign sig_1024 = sig_823 ^ sig_947;
assign sig_1025 = sig_989 | sig_970;
assign sig_1026 = sig_925 ^ sig_838;
assign sig_1027 = sig_920 & sig_714;
assign sig_1028 = sig_945 ^ sig_687;
assign sig_1029 = sig_871 & sig_1014;
assign sig_1030 = sig_936 ^ sig_878;
assign sig_1032 = sig_67 & sig_988;
assign sig_1033 = sig_961 ^ sig_735;
assign sig_1034 = sig_953 ^ sig_841;
assign sig_1036 = sig_953 | sig_841;
assign sig_1037 = sig_876 & sig_1024;
assign sig_1038 = sig_881 | sig_951;
assign sig_1039 = sig_992 ^ sig_722;
assign sig_1040 = sig_943 ^ sig_120;
assign sig_1041 = sig_950 ^ sig_949;
assign sig_1042 = sig_958 & sig_1022;
assign sig_1045 = sig_934 & sig_1027;
assign sig_1046 = sig_966 ^ sig_636;
assign sig_1047 = sig_998 | sig_960;
assign sig_1049 = sig_983 ^ sig_862;
assign sig_1050 = sig_823 & sig_947;
assign sig_1051 = sig_978 | sig_1009;
assign sig_1053 = sig_959 & sig_975;
assign sig_1054 = sig_969 ^ sig_758;
assign sig_1055 = sig_967 ^ sig_754;
assign sig_1056 = sig_962 & sig_695;
assign sig_1058 = sig_996 ^ sig_909;
assign sig_1059 = sig_972 & sig_515;
assign sig_1060 = sig_1011 | sig_940;
assign sig_1061 = sig_992 & sig_722;
assign sig_1062 = sig_1025 ^ sig_684;
assign sig_1063 = sig_985 ^ sig_764;
assign sig_1065 = sig_961 & sig_735;
assign sig_1066 = sig_839 | sig_991;
assign sig_1068 = sig_1025 & sig_684;
assign sig_1069 = sig_988 ^ sig_67;
assign sig_1070 = sig_972 ^ sig_515;
assign sig_1072 = sig_1007 ^ sig_794;
assign sig_1073 = sig_918 & sig_1041;
assign sig_1074 = sig_1038 ^ sig_646;
assign sig_1076 = sig_134 & sig_1049;
assign sig_1078 = sig_983 & sig_862;
assign sig_1079 = sig_987 | sig_1004;
assign sig_1080 = sig_1021 | sig_1032;
assign sig_1082 = sig_1024 ^ sig_876;
assign sig_1084 = sig_1020 & sig_405;
assign sig_1085 = sig_1062 ^ sig_99;
assign sig_1086 = sig_1006 ^ sig_98;
assign sig_1087 = sig_180 & sig_1033;
assign sig_1088 = sig_1014 ^ sig_871;
assign sig_1089 = sig_794 & sig_1007;
assign sig_1090 = sig_974 | sig_1073;
assign sig_1091 = sig_99 & sig_1062;
assign sig_1092 = sig_1000 & sig_691;
assign sig_1093 = sig_1056 | sig_1002;
assign sig_1094 = sig_929 & sig_1018;
assign sig_1095 = sig_1047 ^ sig_666;
assign sig_1096 = sig_941 | sig_1012;
assign sig_1098 = sig_161 & sig_1039;
assign sig_1100 = sig_1065 | sig_1087;
assign sig_1102 = sig_928 | sig_1013;
assign sig_1103 = sig_934 ^ sig_1027;
assign sig_1105 = sig_1072 ^ sig_1066;
assign sig_1106 = sig_1047 & sig_666;
assign sig_1107 = sig_1053 | sig_1029;
assign sig_1108 = sig_1020 ^ sig_405;
assign sig_1109 = sig_1028 ^ sig_36;
assign sig_1111 = sig_958 ^ sig_1022;
assign sig_1112 = sig_36 & sig_1028;
assign sig_1113 = sig_337 & sig_1095;
assign sig_1114 = sig_1050 | sig_1037;
assign sig_1115 = sig_1082 & sig_1107;
assign sig_1117 = sig_1105 ^ sig_901;
assign sig_1119 = sig_1033 ^ sig_180;
assign sig_1120 = sig_757 & sig_1034;
assign sig_1121 = sig_96 & sig_1074;
assign sig_1122 = sig_1068 | sig_1091;
assign sig_1123 = sig_1038 & sig_646;
assign sig_1124 = sig_1039 ^ sig_161;
assign sig_1125 = sig_1058 ^ sig_1079;
assign sig_1126 = sig_80 & sig_1108;
assign sig_1127 = sig_1106 | sig_1113;
assign sig_1129 = sig_1103 ^ sig_1086;
assign sig_1130 = sig_1092 | sig_1023;
assign sig_1131 = sig_742 & sig_1094;
assign sig_1132 = sig_956 ^ sig_1051;
assign sig_1133 = sig_956 & sig_1051;
assign sig_1134 = sig_1049 ^ sig_134;
assign sig_1135 = sig_1041 ^ sig_918;
assign sig_1136 = sig_1055 ^ sig_860;
assign sig_1137 = sig_979 & sig_1114;
assign sig_1139 = sig_860 & sig_1055;
assign sig_1140 = sig_1132 ^ sig_1026;
assign sig_1141 = sig_1058 & sig_1079;
assign sig_1142 = sig_1060 ^ sig_702;
assign sig_1145 = sig_1093 & sig_354;
assign sig_1146 = sig_1123 | sig_1121;
assign sig_1147 = sig_927 & sig_1102;
assign sig_1148 = sig_206 & sig_1070;
assign sig_1149 = sig_1060 & sig_702;
assign sig_1150 = sig_1078 | sig_1076;
assign sig_1151 = sig_1072 & sig_1066;
assign sig_1152 = sig_1074 ^ sig_96;
assign sig_1153 = sig_1084 | sig_1126;
assign sig_1154 = sig_1070 ^ sig_206;
assign sig_1155 = sig_1026 & sig_1132;
assign sig_1156 = sig_1142 ^ sig_285;
assign sig_1158 = sig_957 | sig_1089;
assign sig_1159 = sig_1017 & sig_1125;
assign sig_1160 = sig_1125 ^ sig_1017;
assign sig_1161 = sig_1093 ^ sig_354;
assign sig_1162 = sig_383 ^ sig_1154;
assign sig_1163 = sig_214 & sig_1094;
assign sig_1164 = sig_1095 ^ sig_337;
assign sig_1165 = sig_1133 | sig_1155;
assign sig_1166 = sig_1040 & sig_1111;
assign sig_1167 = sig_901 & sig_1105;
assign sig_1169 = sig_1061 | sig_1098;
assign sig_1170 = sig_1141 | sig_1159;
assign sig_1171 = sig_981 ^ sig_1124;
assign sig_1172 = sig_1082 ^ sig_1107;
assign sig_1174 = sig_1108 ^ sig_80;
assign sig_1175 = sig_1134 & sig_1054;
assign sig_1176 = sig_285 & sig_1142;
assign sig_1177 = sig_927 ^ sig_1102;
assign sig_1178 = sig_1135 ^ sig_1165;
assign sig_1180 = sig_1036 | sig_1120;
assign sig_1181 = sig_965 ^ sig_1119;
assign sig_1182 = sig_1046 & sig_1172;
assign sig_1183 = sig_1042 | sig_1166;
assign sig_1185 = sig_1140 & sig_1170;
assign sig_1186 = sig_979 ^ sig_1114;
assign sig_1187 = sig_1140 ^ sig_1170;
assign sig_1188 = sig_1086 & sig_1103;
assign sig_1189 = sig_1172 ^ sig_1046;
assign sig_1190 = sig_1111 ^ sig_1040;
assign sig_1191 = sig_1151 | sig_1167;
assign sig_1192 = sig_1005 | sig_1112;
assign sig_1193 = sig_1178 ^ sig_1156;
assign sig_1194 = sig_1135 & sig_1165;
assign sig_1195 = sig_971 | sig_1139;
assign sig_1196 = sig_1119 & sig_965;
assign sig_1197 = sig_1149 | sig_1176;
assign sig_1199 = sig_1054 ^ sig_1134;
assign sig_1200 = sig_1063 ^ sig_1158;
assign sig_1201 = sig_1124 & sig_981;
assign sig_1202 = sig_541 & sig_1163;
assign sig_1203 = sig_1136 & sig_942;
assign sig_1204 = sig_1195 ^ sig_656;
assign sig_1205 = sig_1154 & sig_383;
assign sig_1206 = sig_1177 ^ sig_1174;
assign sig_1207 = sig_1115 | sig_1182;
assign sig_1209 = sig_942 ^ sig_1136;
assign sig_1210 = sig_1088 & sig_1180;
assign sig_1213 = sig_1131 | sig_1202;
assign sig_1214 = sig_1199 ^ sig_1183;
assign sig_1215 = sig_1174 & sig_1177;
assign sig_1216 = sig_919 | sig_1203;
assign sig_1218 = sig_1162 & sig_1196;
assign sig_1219 = sig_1181 ^ sig_1201;
assign sig_1220 = sig_718 & sig_1205;
assign sig_1221 = sig_1059 | sig_1148;
assign sig_1222 = sig_718 ^ sig_1205;
assign sig_1223 = sig_1063 & sig_1158;
assign sig_1225 = sig_1162 ^ sig_1196;
assign sig_1226 = sig_1171 ^ sig_1175;
assign sig_1227 = sig_1030 & sig_1216;
assign sig_1231 = sig_532 & sig_930;
assign sig_1232 = sig_1209 & sig_1090;
assign sig_1233 = sig_1222 ^ sig_1221;
assign sig_1234 = sig_907 & sig_1200;
assign sig_1235 = sig_1186 ^ sig_980;
assign sig_1237 = sig_1225 ^ sig_1100;
assign sig_1238 = sig_1199 & sig_1183;
assign sig_1240 = sig_1045 | sig_1188;
assign sig_1242 = sig_980 & sig_1186;
assign sig_1244 = sig_1200 ^ sig_907;
assign sig_1245 = sig_1209 ^ sig_1090;
assign sig_1246 = sig_1169 & sig_1219;
assign sig_1247 = sig_1214 ^ sig_1010;
assign sig_1248 = sig_1156 & sig_1178;
assign sig_1250 = sig_1171 & sig_1175;
assign sig_1251 = sig_1223 | sig_1234;
assign sig_1252 = sig_1187 ^ sig_1085;
assign sig_1253 = sig_1235 & sig_1207;
assign sig_1254 = sig_1147 | sig_1215;
assign sig_1256 = sig_1088 ^ sig_1180;
assign sig_1258 = sig_1150 & sig_1226;
assign sig_1259 = sig_1085 & sig_1187;
assign sig_1260 = sig_1235 ^ sig_1207;
assign sig_1262 = sig_1030 ^ sig_1216;
assign sig_1264 = sig_1181 & sig_1201;
assign sig_1266 = sig_1160 ^ sig_1251;
assign sig_1267 = sig_995 & sig_1256;
assign sig_1268 = sig_1010 & sig_1214;
assign sig_1269 = sig_1219 ^ sig_1169;
assign sig_1270 = sig_1069 & sig_1266;
assign sig_1271 = sig_1137 | sig_1242;
assign sig_1272 = sig_50 & sig_1204;
assign sig_1273 = sig_1226 ^ sig_1150;
assign sig_1274 = sig_1244 ^ sig_1191;
assign sig_1275 = sig_1204 ^ sig_50;
assign sig_1277 = sig_1195 & sig_656;
assign sig_1280 = sig_1256 ^ sig_995;
assign sig_1281 = sig_1238 | sig_1268;
assign sig_1282 = sig_1210 | sig_1267;
assign sig_1283 = sig_1161 & sig_1260;
assign sig_1284 = sig_1109 & sig_1245;
assign sig_1285 = sig_1129 & sig_1254;
assign sig_1286 = sig_1129 ^ sig_1254;
assign sig_1287 = sig_1286 ^ sig_1153;
assign sig_1288 = sig_1221 & sig_1222;
assign sig_1289 = sig_1253 | sig_1283;
assign sig_1290 = sig_1264 | sig_1246;
assign sig_1291 = sig_1277 | sig_1272;
assign sig_1292 = sig_1220 | sig_1288;
assign sig_1293 = sig_1100 & sig_1225;
assign sig_1295 = sig_1245 ^ sig_1109;
assign sig_1296 = sig_1218 | sig_1293;
assign sig_1297 = sig_1250 | sig_1258;
assign sig_1299 = sig_1273 & sig_1281;
assign sig_1300 = sig_1015 & sig_649;
assign sig_1301 = sig_1262 ^ sig_1275;
assign sig_1302 = sig_1190 ^ sig_1240;
assign sig_1303 = sig_900 & sig_1213;
assign sig_1304 = sig_1189 & sig_1282;
assign sig_1305 = sig_1266 ^ sig_1069;
assign sig_1306 = sig_1275 & sig_1262;
assign sig_1307 = sig_1185 | sig_1259;
assign sig_1308 = sig_1130 & sig_1302;
assign sig_1309 = sig_1153 & sig_1286;
assign sig_1310 = sig_1274 ^ sig_1152;
assign sig_1311 = sig_1233 ^ sig_1296;
assign sig_1312 = sig_1194 | sig_1248;
assign sig_1313 = sig_1269 ^ sig_1297;
assign sig_1314 = sig_1237 ^ sig_1290;
assign sig_1316 = sig_1273 ^ sig_1281;
assign sig_1317 = sig_1227 | sig_1306;
assign sig_1318 = sig_1189 ^ sig_1282;
assign sig_1319 = sig_1260 ^ sig_1161;
assign sig_1320 = sig_1190 & sig_1240;
assign sig_1321 = sig_1244 & sig_1191;
assign sig_1323 = sig_1232 | sig_1284;
assign sig_1324 = sig_1280 | sig_1213;
assign sig_1325 = sig_1160 & sig_1251;
assign sig_1327 = sig_1117 ^ sig_1271;
assign sig_1328 = sig_774 & sig_1292;
assign sig_1329 = sig_1313 & sig_1299;
assign sig_1330 = sig_1028 | sig_1106;
assign sig_1331 = sig_1302 ^ sig_1130;
assign sig_1332 = sig_1117 & sig_1271;
assign sig_1335 = sig_1285 | sig_1309;
assign sig_1337 = sig_1193 ^ sig_1307;
assign sig_1338 = sig_1295 & sig_1312;
assign sig_1339 = sig_1231 & sig_1300;
assign sig_1340 = sig_1152 & sig_1274;
assign sig_1342 = sig_1193 & sig_1307;
assign sig_1343 = sig_1301 & sig_1323;
assign sig_1344 = sig_1301 ^ sig_1323;
assign sig_1345 = sig_1344 ^ sig_1192;
assign sig_1346 = sig_1164 & sig_1327;
assign sig_1347 = sig_1295 ^ sig_1312;
assign sig_1349 = sig_1233 & sig_1296;
assign sig_1350 = sig_1206 & sig_1317;
assign sig_1351 = sig_774 ^ sig_1292;
assign sig_1352 = sig_1347 ^ sig_1197;
assign sig_1353 = sig_1313 & sig_1316;
assign sig_1354 = sig_1337 ^ sig_1122;
assign sig_1355 = sig_1320 | sig_1308;
assign sig_1356 = sig_1318 ^ sig_1096;
assign sig_1357 = sig_1237 & sig_1290;
assign sig_1359 = sig_1096 & sig_1318;
assign sig_1360 = sig_1311 & sig_1314;
assign sig_1361 = sig_1324 ^ sig_994;
assign sig_1362 = sig_1269 & sig_1297;
assign sig_1363 = sig_1206 ^ sig_1317;
assign sig_1364 = sig_928 & sig_1339;
assign sig_1365 = sig_994 & sig_1324;
assign sig_1366 = sig_1332 | sig_1346;
assign sig_1367 = sig_1122 & sig_1337;
assign sig_1368 = sig_1363 ^ sig_1291;
assign sig_1369 = sig_1321 | sig_1340;
assign sig_1370 = sig_1310 & sig_1366;
assign sig_1371 = sig_1247 & sig_1355;
assign sig_1372 = sig_1325 | sig_1270;
assign sig_1374 = sig_1331 & sig_1335;
assign sig_1377 = sig_1291 & sig_1363;
assign sig_1379 = sig_1327 ^ sig_1164;
assign sig_1380 = sig_1192 & sig_1344;
assign sig_1382 = sig_1379 ^ sig_1289;
assign sig_1383 = sig_1247 ^ sig_1355;
assign sig_1384 = sig_1197 & sig_1347;
assign sig_1385 = sig_1383 & sig_1374;
assign sig_1386 = sig_1310 ^ sig_1366;
assign sig_1387 = sig_1342 | sig_1367;
assign sig_1388 = sig_1331 ^ sig_1335;
assign sig_1389 = sig_1361 | sig_1339;
assign sig_1390 = sig_1343 | sig_1380;
assign sig_1391 = sig_1305 ^ sig_1369;
assign sig_1393 = sig_1311 & sig_1357;
assign sig_1394 = sig_1252 ^ sig_1372;
assign sig_1395 = sig_1368 ^ sig_1390;
assign sig_1397 = sig_1338 | sig_1384;
assign sig_1398 = sig_1362 | sig_1329;
assign sig_1400 = sig_1345 ^ sig_1397;
assign sig_1401 = sig_1352 ^ sig_1387;
assign sig_1402 = sig_1350 | sig_1377;
assign sig_1403 = sig_1252 & sig_1372;
assign sig_1404 = sig_1303 | sig_1365;
assign sig_1405 = sig_1394 ^ sig_1080;
assign sig_1406 = sig_1400 & sig_1401;
assign sig_1407 = sig_1371 | sig_1385;
assign sig_1408 = sig_1304 | sig_1359;
assign sig_1409 = sig_1379 & sig_1289;
assign sig_1410 = sig_1080 & sig_1394;
assign sig_1411 = sig_1127 & sig_1386;
assign sig_1412 = sig_1383 & sig_1388;
assign sig_1413 = sig_1353 & sig_1412;
assign sig_1414 = sig_1146 & sig_1391;
assign sig_1415 = sig_1305 & sig_1369;
assign sig_1416 = sig_1356 & sig_1404;
assign sig_1417 = sig_1319 ^ sig_1408;
assign sig_1419 = sig_1319 & sig_1408;
assign sig_1421 = sig_1382 ^ sig_1145;
assign sig_1422 = sig_1145 & sig_1382;
assign sig_1423 = sig_1409 | sig_1422;
assign sig_1424 = sig_1386 ^ sig_1127;
assign sig_1425 = sig_1424 & sig_1423;
assign sig_1427 = sig_1287 & sig_1402;
assign sig_1428 = sig_1370 | sig_1411;
assign sig_1429 = sig_1391 ^ sig_1146;
assign sig_1430 = sig_1353 & sig_1407;
assign sig_1431 = sig_1368 & sig_1390;
assign sig_1432 = sig_1415 | sig_1414;
assign sig_1433 = sig_1429 & sig_1428;
assign sig_1435 = sig_1345 & sig_1397;
assign sig_1436 = sig_1417 & sig_1416;
assign sig_1437 = sig_1403 | sig_1410;
assign sig_1438 = sig_1352 & sig_1387;
assign sig_1439 = sig_1421 & sig_1419;
assign sig_1440 = sig_1349 | sig_1393;
assign sig_1441 = sig_1287 ^ sig_1402;
assign sig_1442 = sig_1356 ^ sig_1404;
assign sig_1443 = sig_1442 | sig_1364;
assign sig_1444 = sig_1398 | sig_1430;
assign sig_1447 = sig_1405 & sig_1432;
assign sig_1449 = sig_1354 & sig_1437;
assign sig_1450 = sig_1400 & sig_1438;
assign sig_1451 = sig_1424 ^ sig_1423;
assign sig_1452 = sig_1441 & sig_1431;
assign sig_1454 = sig_1429 ^ sig_1428;
assign sig_1455 = sig_401 & sig_1202;
assign sig_1456 = sig_1417 ^ sig_1416;
assign sig_1457 = sig_333 & sig_1094;
assign sig_1458 = sig_897 & sig_1457;
assign sig_1459 = sig_1421 ^ sig_1419;
assign sig_1461 = sig_1459 & sig_1436;
assign sig_1462 = sig_1405 ^ sig_1432;
assign sig_1464 = sig_1454 & sig_1425;
assign sig_1465 = sig_1354 ^ sig_1437;
assign sig_1467 = sig_1465 & sig_1447;
assign sig_1468 = sig_1441 & sig_1395;
assign sig_1469 = sig_1459 & sig_1456;
assign sig_1471 = sig_1389 | sig_1455;
assign sig_1472 = sig_1465 & sig_1462;
assign sig_1473 = sig_1427 | sig_1452;
assign sig_1474 = sig_1454 & sig_1451;
assign sig_1475 = sig_1435 | sig_1450;
assign sig_1477 = sig_1472 & sig_1474;
assign sig_1478 = sig_1468 & sig_1406;
assign sig_1479 = sig_1439 | sig_1461;
assign sig_1481 = sig_813 & sig_1458;
assign sig_1483 = sig_1449 | sig_1467;
assign sig_1484 = sig_1478 & sig_1477;
assign sig_1485 = sig_1433 | sig_1464;
assign sig_1489 = sig_1472 & sig_1485;
assign sig_1490 = sig_1483 | sig_1489;
assign sig_1491 = sig_1468 & sig_1475;
assign sig_1492 = sig_1443 & sig_1471;
assign sig_1493 = sig_1473 | sig_1491;
assign sig_1497 = sig_1469 & sig_1492;
assign sig_1498 = A[10] & sig_146;
assign sig_1499 = sig_1479 | sig_1461;
assign sig_1500 = sig_1497 & sig_1498;
assign sig_1501 = sig_1478 & sig_1490;
assign sig_1502 = sig_1493 | sig_1501;
assign sig_1503 = sig_1498 & sig_1330;
assign sig_1504 = sig_1500 & sig_1330;
assign sig_1505 = sig_1127 | sig_580;
assign sig_1506 = sig_1505 | sig_1503;
assign sig_1507 = sig_1471 ^ sig_1506;
assign sig_1508 = sig_1471 & sig_1506;
assign sig_1509 = sig_1497 & sig_1505;
assign sig_1510 = sig_1492 & sig_1506;
assign sig_1511 = sig_1481 | sig_1510;
assign sig_1512 = sig_1457 | sig_1508;
assign sig_1513 = sig_1456 & sig_1511;
assign sig_1514 = sig_1499 | sig_1509;
assign sig_1515 = sig_1443 ^ sig_1512;
assign sig_1516 = sig_1456 ^ sig_1511;
assign sig_1517 = sig_1514 | sig_1504;
assign sig_1518 = sig_1436 ^ sig_1513;
assign sig_1519 = sig_1451 & sig_1517;
assign sig_1520 = sig_1484 & sig_1517;
assign sig_1521 = sig_1477 & sig_1517;
assign sig_1522 = sig_1451 ^ sig_1517;
assign sig_1523 = sig_1490 | sig_1521;
assign sig_1524 = sig_1406 & sig_1523;
assign sig_1525 = sig_1474 & sig_1517;
assign sig_1526 = sig_1459 ^ sig_1518;
assign sig_1527 = sig_1425 | sig_1519;
assign sig_1528 = sig_1502 | sig_1520;
assign sig_1529 = sig_1475 | sig_1524;
assign sig_1530 = sig_1401 & sig_1523;
assign sig_1531 = sig_1412 & sig_1528;
assign sig_1532 = sig_1395 & sig_1529;
assign sig_1533 = sig_1388 ^ sig_1528;
assign sig_1534 = sig_1407 | sig_1531;
assign sig_1535 = sig_1395 ^ sig_1529;
assign sig_1536 = sig_1485 | sig_1525;
assign sig_1537 = sig_1401 ^ sig_1523;
assign sig_1538 = sig_1388 & sig_1528;
assign sig_1539 = sig_1413 & sig_1528;
assign sig_1540 = sig_1316 & sig_1534;
assign sig_1541 = sig_1454 ^ sig_1527;
assign sig_1542 = sig_1431 | sig_1532;
assign sig_1543 = sig_1462 ^ sig_1536;
assign sig_1544 = sig_1438 | sig_1530;
assign sig_1545 = sig_1299 | sig_1540;
assign sig_1546 = sig_1316 ^ sig_1534;
assign sig_1547 = sig_1444 | sig_1539;
assign sig_1548 = sig_1374 | sig_1538;
assign sig_1549 = sig_1441 ^ sig_1542;
assign sig_1550 = sig_1462 & sig_1536;
assign sig_1551 = sig_1314 & sig_1547;
assign sig_1552 = sig_1400 ^ sig_1544;
assign sig_1553 = sig_1357 | sig_1551;
assign sig_1554 = sig_1447 | sig_1550;
assign sig_1555 = sig_1465 ^ sig_1554;
assign sig_1556 = sig_1313 ^ sig_1545;
assign sig_1557 = sig_1311 ^ sig_1553;
assign sig_1558 = sig_1314 ^ sig_1547;
assign sig_1559 = sig_1360 & sig_1547;
assign sig_1560 = sig_1383 ^ sig_1548;
assign sig_1561 = sig_1440 | sig_1559;
assign sig_1562 = sig_1351 ^ sig_1561;
assign sig_1563 = sig_1351 & sig_1561;
assign sig_1564 = sig_1328 | sig_1563;
assign sig_1565 = sig_890 | sig_1564;

assign Z[0] = sig_328;
assign Z[1] = sig_802;
assign Z[2] = sig_1511;
assign Z[3] = sig_784;
assign Z[4] = sig_594;
assign Z[5] = sig_1309;
assign Z[6] = sig_748;
assign Z[7] = sig_670;
assign Z[8] = sig_765;
assign Z[9] = sig_852;
assign Z[10] = A[5];
assign Z[11] = sig_168;
assign Z[12] = sig_1507;
assign Z[13] = sig_1515;
assign Z[14] = sig_1516;
assign Z[15] = sig_1526;
assign Z[16] = sig_1522;
assign Z[17] = sig_1541;
assign Z[18] = sig_1543;
assign Z[19] = sig_1555;
assign Z[20] = sig_1537;
assign Z[21] = sig_1552;
assign Z[22] = sig_1535;
assign Z[23] = sig_1549;
assign Z[24] = sig_1533;
assign Z[25] = sig_1560;
assign Z[26] = sig_1546;
assign Z[27] = sig_1556;
assign Z[28] = sig_1558;
assign Z[29] = sig_1557;
assign Z[30] = sig_1562;
assign Z[31] = sig_1565;

endmodule



